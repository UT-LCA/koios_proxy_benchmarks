
module top (input clk, input reset,input [602:0] top_inp, output [419:0] top_outp); 
 


 wire [251:0] inp_fifo1;
wire [247:0] outp_fifo1;

fifo_512_60bit_module_4 fifo1 (.clk(clk),.reset(reset),.inp(inp_fifo1),.outp(outp_fifo1)); 


 wire [85:0] inp_fifo2;
wire [83:0] outp_fifo2;

fifo_256_40bit_module_2 fifo2 (.clk(clk),.reset(reset),.inp(inp_fifo2),.outp(outp_fifo2)); 


 wire [1059:0] inp_dot1;
wire [1003:0] outp_dot1;

tensor_block_int8_module_4 dot1 (.clk(clk),.reset(reset),.inp(inp_dot1),.outp(outp_dot1)); 
wire [331:0] inp_interface_2; 
wire [1059:0] outp_interface_2; 

interface_2 inst_interface_2(.clk(clk),.reset(reset),.inp(inp_interface_2),.outp(outp_interface_2)); 


 wire [2119:0] inp_dot2;
wire [2007:0] outp_dot2;

tensor_block_int8_module_8 dot2 (.clk(clk),.reset(reset),.inp(inp_dot2),.outp(outp_dot2)); 
wire [2315:0] inp_interface_3; 
wire [2119:0] outp_interface_3; 

interface_3 inst_interface_3(.clk(clk),.reset(reset),.inp(inp_interface_3),.outp(outp_interface_3)); 


 wire [1775:0] inp_dspch1;
wire [221:0] outp_dspch1;

dsp_chain_4_int_sop_2_module_6 dspch1 (.clk(clk),.reset(reset),.inp(inp_dspch1),.outp(outp_dspch1)); 
wire [331:0] inp_interface_4; 
wire [1775:0] outp_interface_4; 

interface_4 inst_interface_4(.clk(clk),.reset(reset),.inp(inp_interface_4),.outp(outp_interface_4)); 


 wire [1031:0] inp_fifo3;
wire [1007:0] outp_fifo3;

fifo_256_40bit_module_24 fifo3 (.clk(clk),.reset(reset),.inp(inp_fifo3),.outp(outp_fifo3)); 
wire [1003:0] inp_interface_5; 
wire [1031:0] outp_interface_5; 

interface_5 inst_interface_5(.clk(clk),.reset(reset),.inp(inp_interface_5),.outp(outp_interface_5)); 


 wire [2519:0] inp_fifo4;
wire [2479:0] outp_fifo4;

fifo_512_60bit_module_40 fifo4 (.clk(clk),.reset(reset),.inp(inp_fifo4),.outp(outp_fifo4)); 
wire [1003:0] inp_interface_6; 
wire [2519:0] outp_interface_6; 

interface_6 inst_interface_6(.clk(clk),.reset(reset),.inp(inp_interface_6),.outp(outp_interface_6)); 


 wire [1133:0] inp_fifo5;
wire [1115:0] outp_fifo5;

fifo_256_60bit_module_18 fifo5 (.clk(clk),.reset(reset),.inp(inp_fifo5),.outp(outp_fifo5)); 
wire [2007:0] inp_interface_7; 
wire [1133:0] outp_interface_7; 

interface_7 inst_interface_7(.clk(clk),.reset(reset),.inp(inp_interface_7),.outp(outp_interface_7)); 


 wire [1117:0] inp_fifo6;
wire [1091:0] outp_fifo6;

fifo_512_40bit_module_26 fifo6 (.clk(clk),.reset(reset),.inp(inp_fifo6),.outp(outp_fifo6)); 
wire [2007:0] inp_interface_8; 
wire [1117:0] outp_interface_8; 

interface_8 inst_interface_8(.clk(clk),.reset(reset),.inp(inp_interface_8),.outp(outp_interface_8)); 


 wire [3551:0] inp_dspch4;
wire [591:0] outp_dspch4;

dsp_chain_3_int_sop_2_module_16 dspch4 (.clk(clk),.reset(reset),.inp(inp_dspch4),.outp(outp_dspch4)); 
wire [1007:0] inp_interface_9; 
wire [3551:0] outp_interface_9; 

interface_9 inst_interface_9(.clk(clk),.reset(reset),.inp(inp_interface_9),.outp(outp_interface_9)); 


 wire [1059:0] inp_dot3;
wire [1003:0] outp_dot3;

tensor_block_int8_module_4 dot3 (.clk(clk),.reset(reset),.inp(inp_dot3),.outp(outp_dot3)); 
wire [2479:0] inp_interface_10; 
wire [1059:0] outp_interface_10; 

interface_10 inst_interface_10(.clk(clk),.reset(reset),.inp(inp_interface_10),.outp(outp_interface_10)); 


 wire [171:0] inp_fifo8;
wire [167:0] outp_fifo8;

fifo_256_40bit_module_4 fifo8 (.clk(clk),.reset(reset),.inp(inp_fifo8),.outp(outp_fifo8)); 
wire [1595:0] inp_interface_11; 
wire [171:0] outp_interface_11; 

interface_11 inst_interface_11(.clk(clk),.reset(reset),.inp(inp_interface_11),.outp(outp_interface_11)); 


 wire [2367:0] inp_dspch3;
wire [295:0] outp_dspch3;

dsp_chain_4_int_sop_2_module_8 dspch3 (.clk(clk),.reset(reset),.inp(inp_dspch3),.outp(outp_dspch3)); 
wire [2207:0] inp_interface_12; 
wire [2367:0] outp_interface_12; 

interface_12 inst_interface_12(.clk(clk),.reset(reset),.inp(inp_interface_12),.outp(outp_interface_12)); 


 wire [264:0] inp_dot4;
wire [250:0] outp_dot4;

tensor_block_int8_module_1 dot4 (.clk(clk),.reset(reset),.inp(inp_dot4),.outp(outp_dot4)); 


 wire [2015:0] inp_fifo7;
wire [1983:0] outp_fifo7;

fifo_512_60bit_module_32 fifo7 (.clk(clk),.reset(reset),.inp(inp_fifo7),.outp(outp_fifo7)); 
wire [250:0] inp_interface_14; 
wire [2015:0] outp_interface_14; 

interface_14 inst_interface_14(.clk(clk),.reset(reset),.inp(inp_interface_14),.outp(outp_interface_14)); 


 wire [3699:0] inp_dspch2;
wire [924:0] outp_dspch2;

dsp_chain_2_int_sop_2_module_25 dspch2 (.clk(clk),.reset(reset),.inp(inp_dspch2),.outp(outp_dspch2)); 
wire [3075:0] inp_interface_15; 
wire [3699:0] outp_interface_15; 

interface_15 inst_interface_15(.clk(clk),.reset(reset),.inp(inp_interface_15),.outp(outp_interface_15)); 


 wire [257:0] inp_fifo9;
wire [251:0] outp_fifo9;

fifo_256_40bit_module_6 fifo9 (.clk(clk),.reset(reset),.inp(inp_fifo9),.outp(outp_fifo9)); 
wire [1220:0] inp_interface_16; 
wire [257:0] outp_interface_16; 

interface_16 inst_interface_16(.clk(clk),.reset(reset),.inp(inp_interface_16),.outp(outp_interface_16)); 

assign inp_fifo1 = top_inp[251:0]; 

assign inp_fifo2 = top_inp[337:252]; 

assign inp_dot1 = outp_interface_2; 
assign inp_interface_2 = {outp_fifo1,outp_fifo2}; 
 

assign inp_dot2 = outp_interface_3; 
assign inp_interface_3 = {outp_fifo1,outp_fifo2,outp_fifo7}; 
 

assign inp_dspch1 = outp_interface_4; 
assign inp_interface_4 = {outp_fifo1,outp_fifo2}; 
 

assign inp_fifo3 = outp_interface_5; 
assign inp_interface_5 = {outp_dot1}; 
 

assign inp_fifo4 = outp_interface_6; 
assign inp_interface_6 = {outp_dot1}; 
 

assign inp_fifo5 = outp_interface_7; 
assign inp_interface_7 = {outp_dot2}; 
 

assign inp_fifo6 = outp_interface_8; 
assign inp_interface_8 = {outp_dot2}; 
 

assign inp_dspch4 = outp_interface_9; 
assign inp_interface_9 = {outp_fifo3}; 
 

assign inp_dot3 = outp_interface_10; 
assign inp_interface_10 = {outp_fifo4}; 
 

assign inp_fifo8 = outp_interface_11; 
assign top_outp[167:0] = outp_fifo8; 
assign inp_interface_11 = {outp_dspch4,outp_dot3}; 
 

assign inp_dspch3 = outp_interface_12; 
assign inp_interface_12 = {outp_fifo5,outp_fifo6}; 
 

assign inp_dot4 = top_inp[602:338]; 

assign inp_fifo7 = outp_interface_14; 
assign inp_interface_14 = {outp_dot4}; 
 

assign inp_dspch2 = outp_interface_15; 
assign inp_interface_15 = {outp_fifo7,outp_fifo6}; 
 

assign inp_fifo9 = outp_interface_16; 
assign top_outp[419:168] = outp_fifo9; 
assign inp_interface_16 = {outp_dspch2,outp_dspch3}; 
 

 endmodule 


module interface_2(input [331:0] inp, output reg [1059:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[331:0] <= inp ; 
outp[663:332] <= inp ; 
outp[995:664] <= inp ; 
outp[1059:996] <= inp[63:0] ; 
end 
endmodule 

module interface_3(input [2315:0] inp, output reg [2119:0] outp, input clk, input reset);
reg [2315:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1157:0]intermediate_reg_1; 
 
fsm fsm_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
fsm fsm_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156])); 
xor_module xor_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155])); 
fsm fsm_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154])); 
fsm fsm_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153])); 
fsm fsm_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152])); 
fsm fsm_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147])); 
xor_module xor_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146])); 
fsm fsm_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145])); 
fsm fsm_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143])); 
fsm fsm_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140])); 
fsm fsm_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139])); 
fsm fsm_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137])); 
fsm fsm_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136])); 
fsm fsm_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133])); 
xor_module xor_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132])); 
fsm fsm_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
fsm fsm_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129])); 
fsm fsm_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128])); 
fsm fsm_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127])); 
fsm fsm_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126])); 
fsm fsm_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
fsm fsm_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122])); 
fsm fsm_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120])); 
fsm fsm_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
fsm fsm_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115])); 
fsm fsm_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113])); 
fsm fsm_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111])); 
fsm fsm_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110])); 
fsm fsm_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109])); 
fsm fsm_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
xor_module xor_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106])); 
xor_module xor_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
fsm fsm_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
fsm fsm_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
fsm fsm_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
fsm fsm_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100])); 
fsm fsm_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097])); 
fsm fsm_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096])); 
xor_module xor_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095])); 
fsm fsm_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
fsm fsm_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
fsm fsm_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090])); 
xor_module xor_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088])); 
fsm fsm_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
fsm fsm_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086])); 
xor_module xor_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085])); 
fsm fsm_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084])); 
xor_module xor_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
fsm fsm_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082])); 
fsm fsm_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081])); 
fsm fsm_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080])); 
xor_module xor_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
fsm fsm_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076])); 
fsm fsm_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075])); 
fsm fsm_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069])); 
fsm fsm_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066])); 
fsm fsm_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063])); 
xor_module xor_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061])); 
fsm fsm_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060])); 
fsm fsm_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059])); 
fsm fsm_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055])); 
xor_module xor_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054])); 
xor_module xor_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051])); 
fsm fsm_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
fsm fsm_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046])); 
xor_module xor_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
xor_module xor_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
fsm fsm_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
fsm fsm_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041])); 
fsm fsm_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039])); 
xor_module xor_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038])); 
fsm fsm_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036])); 
fsm fsm_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035])); 
fsm fsm_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033])); 
fsm fsm_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032])); 
fsm fsm_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
fsm fsm_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030])); 
xor_module xor_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026])); 
fsm fsm_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024])); 
xor_module xor_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
fsm fsm_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022])); 
xor_module xor_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021])); 
fsm fsm_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
fsm fsm_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017])); 
fsm fsm_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
xor_module xor_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
xor_module xor_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013])); 
fsm fsm_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011])); 
fsm fsm_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010])); 
xor_module xor_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009])); 
fsm fsm_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006])); 
fsm fsm_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
fsm fsm_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
xor_module xor_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
fsm fsm_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991])); 
fsm fsm_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
xor_module xor_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
fsm fsm_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
fsm fsm_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
fsm fsm_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
fsm fsm_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
xor_module xor_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
xor_module xor_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
fsm fsm_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
fsm fsm_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975])); 
xor_module xor_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974])); 
fsm fsm_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
xor_module xor_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
xor_module xor_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971])); 
fsm fsm_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
xor_module xor_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
xor_module xor_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
fsm fsm_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
fsm fsm_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
xor_module xor_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
xor_module xor_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959])); 
fsm fsm_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
fsm fsm_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954])); 
fsm fsm_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
fsm fsm_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
xor_module xor_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950])); 
fsm fsm_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
xor_module xor_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948])); 
fsm fsm_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
fsm fsm_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
xor_module xor_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
xor_module xor_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
xor_module xor_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
fsm fsm_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
xor_module xor_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
fsm fsm_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
xor_module xor_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
fsm fsm_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
fsm fsm_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
fsm fsm_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
xor_module xor_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
fsm fsm_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
fsm fsm_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
fsm fsm_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
xor_module xor_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
fsm fsm_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
xor_module xor_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
fsm fsm_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
fsm fsm_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
xor_module xor_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
fsm fsm_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
fsm fsm_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
xor_module xor_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
fsm fsm_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
fsm fsm_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
xor_module xor_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
fsm fsm_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
fsm fsm_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
xor_module xor_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
xor_module xor_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
fsm fsm_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
fsm fsm_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
fsm fsm_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
fsm fsm_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
fsm fsm_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
fsm fsm_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
xor_module xor_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886])); 
fsm fsm_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884])); 
xor_module xor_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
xor_module xor_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
fsm fsm_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
fsm fsm_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879])); 
fsm fsm_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
xor_module xor_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
fsm fsm_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
fsm fsm_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
fsm fsm_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
fsm fsm_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
fsm fsm_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
fsm fsm_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
xor_module xor_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
fsm fsm_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
fsm fsm_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865])); 
xor_module xor_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
fsm fsm_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
xor_module xor_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
xor_module xor_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
xor_module xor_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
xor_module xor_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
fsm fsm_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
fsm fsm_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
xor_module xor_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
fsm fsm_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
fsm fsm_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842])); 
fsm fsm_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
xor_module xor_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
fsm fsm_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
fsm fsm_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
xor_module xor_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
xor_module xor_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
fsm fsm_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
fsm fsm_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
fsm fsm_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831])); 
xor_module xor_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
fsm fsm_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
xor_module xor_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
xor_module xor_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
fsm fsm_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823])); 
xor_module xor_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
fsm fsm_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
xor_module xor_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
xor_module xor_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
fsm fsm_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810])); 
xor_module xor_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
xor_module xor_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
fsm fsm_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
fsm fsm_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
fsm fsm_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
xor_module xor_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
fsm fsm_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
fsm fsm_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
xor_module xor_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
fsm fsm_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
xor_module xor_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
fsm fsm_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
xor_module xor_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
xor_module xor_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
xor_module xor_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
fsm fsm_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
xor_module xor_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
fsm fsm_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
fsm fsm_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
fsm fsm_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
xor_module xor_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
fsm fsm_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
fsm fsm_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
xor_module xor_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
fsm fsm_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
fsm fsm_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
xor_module xor_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
xor_module xor_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
fsm fsm_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
fsm fsm_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
xor_module xor_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
fsm fsm_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
xor_module xor_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
xor_module xor_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
xor_module xor_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
fsm fsm_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
xor_module xor_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
xor_module xor_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
xor_module xor_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
fsm fsm_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
xor_module xor_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
xor_module xor_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
xor_module xor_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
xor_module xor_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
fsm fsm_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
xor_module xor_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
xor_module xor_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
xor_module xor_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
fsm fsm_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
fsm fsm_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
fsm fsm_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
fsm fsm_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
fsm fsm_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
fsm fsm_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
fsm fsm_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
fsm fsm_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
fsm fsm_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
fsm fsm_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
fsm fsm_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
xor_module xor_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
fsm fsm_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
fsm fsm_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
fsm fsm_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
xor_module xor_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
fsm fsm_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687])); 
xor_module xor_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
xor_module xor_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
fsm fsm_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
fsm fsm_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
fsm fsm_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
fsm fsm_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
fsm fsm_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
fsm fsm_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
xor_module xor_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
xor_module xor_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
fsm fsm_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
fsm fsm_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
fsm fsm_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
xor_module xor_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
fsm fsm_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
fsm fsm_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
xor_module xor_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
xor_module xor_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
fsm fsm_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
xor_module xor_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
fsm fsm_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
xor_module xor_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
xor_module xor_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
fsm fsm_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
fsm fsm_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
xor_module xor_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
fsm fsm_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
fsm fsm_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
fsm fsm_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
fsm fsm_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640])); 
fsm fsm_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
xor_module xor_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
xor_module xor_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
xor_module xor_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
fsm fsm_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
fsm fsm_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
xor_module xor_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
fsm fsm_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
fsm fsm_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
fsm fsm_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
fsm fsm_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
fsm fsm_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
fsm fsm_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
fsm fsm_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
fsm fsm_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
xor_module xor_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
fsm fsm_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
xor_module xor_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
fsm fsm_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
xor_module xor_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
xor_module xor_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
fsm fsm_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
fsm fsm_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
xor_module xor_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
fsm fsm_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
xor_module xor_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
fsm fsm_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
xor_module xor_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
xor_module xor_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
fsm fsm_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
fsm fsm_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
fsm fsm_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
xor_module xor_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
fsm fsm_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
fsm fsm_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
xor_module xor_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
fsm fsm_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
fsm fsm_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
fsm fsm_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
xor_module xor_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
fsm fsm_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
fsm fsm_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
xor_module xor_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
xor_module xor_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
fsm fsm_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
fsm fsm_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
fsm fsm_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
fsm fsm_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
fsm fsm_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
fsm fsm_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
xor_module xor_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
xor_module xor_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
xor_module xor_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
xor_module xor_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
xor_module xor_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
fsm fsm_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
fsm fsm_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
xor_module xor_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
xor_module xor_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
fsm fsm_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
fsm fsm_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
fsm fsm_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
fsm fsm_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
xor_module xor_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
fsm fsm_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
xor_module xor_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
fsm fsm_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
fsm fsm_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
fsm fsm_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
fsm fsm_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
fsm fsm_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
xor_module xor_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
xor_module xor_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
xor_module xor_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
xor_module xor_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
fsm fsm_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
xor_module xor_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
fsm fsm_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
xor_module xor_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
fsm fsm_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
fsm fsm_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
fsm fsm_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
xor_module xor_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
fsm fsm_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
fsm fsm_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
xor_module xor_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
fsm fsm_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
fsm fsm_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
xor_module xor_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
xor_module xor_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
xor_module xor_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
xor_module xor_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
fsm fsm_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
fsm fsm_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
fsm fsm_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
xor_module xor_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
fsm fsm_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
fsm fsm_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
xor_module xor_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
xor_module xor_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
fsm fsm_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
fsm fsm_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
fsm fsm_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
xor_module xor_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
fsm fsm_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
fsm fsm_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
fsm fsm_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
fsm fsm_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
fsm fsm_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
fsm fsm_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
xor_module xor_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
xor_module xor_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
fsm fsm_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
fsm fsm_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
fsm fsm_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
xor_module xor_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
xor_module xor_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
xor_module xor_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
fsm fsm_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
fsm fsm_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
xor_module xor_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
fsm fsm_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
fsm fsm_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
xor_module xor_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
xor_module xor_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
xor_module xor_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
fsm fsm_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
xor_module xor_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
xor_module xor_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
fsm fsm_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
fsm fsm_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
fsm fsm_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
xor_module xor_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
xor_module xor_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
fsm fsm_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
fsm fsm_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
xor_module xor_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
xor_module xor_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
fsm fsm_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
fsm fsm_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
fsm fsm_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
xor_module xor_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
fsm fsm_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
fsm fsm_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
fsm fsm_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
xor_module xor_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
xor_module xor_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
xor_module xor_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
fsm fsm_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
xor_module xor_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
xor_module xor_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
fsm fsm_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
xor_module xor_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
xor_module xor_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
xor_module xor_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
xor_module xor_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
xor_module xor_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
fsm fsm_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
xor_module xor_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
xor_module xor_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
fsm fsm_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
fsm fsm_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
xor_module xor_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
xor_module xor_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
fsm fsm_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
fsm fsm_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
fsm fsm_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
fsm fsm_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
xor_module xor_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
xor_module xor_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
xor_module xor_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
fsm fsm_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
xor_module xor_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
xor_module xor_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
xor_module xor_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
xor_module xor_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
fsm fsm_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
xor_module xor_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
fsm fsm_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
fsm fsm_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
xor_module xor_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
xor_module xor_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
fsm fsm_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
xor_module xor_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
xor_module xor_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
xor_module xor_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
fsm fsm_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
xor_module xor_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
xor_module xor_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
fsm fsm_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
fsm fsm_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
xor_module xor_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
xor_module xor_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
fsm fsm_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
fsm fsm_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
fsm fsm_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
xor_module xor_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
fsm fsm_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
xor_module xor_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
fsm fsm_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
xor_module xor_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
xor_module xor_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
xor_module xor_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
xor_module xor_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
fsm fsm_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
xor_module xor_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
xor_module xor_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
xor_module xor_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
fsm fsm_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
xor_module xor_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
fsm fsm_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
fsm fsm_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
xor_module xor_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
fsm fsm_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
fsm fsm_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
fsm fsm_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
fsm fsm_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
xor_module xor_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
xor_module xor_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
fsm fsm_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
xor_module xor_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
xor_module xor_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
xor_module xor_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
xor_module xor_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
xor_module xor_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
xor_module xor_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
fsm fsm_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
xor_module xor_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
xor_module xor_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
fsm fsm_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
xor_module xor_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
xor_module xor_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
fsm fsm_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
fsm fsm_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
xor_module xor_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
fsm fsm_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
fsm fsm_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
xor_module xor_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
fsm fsm_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
fsm fsm_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
xor_module xor_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
fsm fsm_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
fsm fsm_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
xor_module xor_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
fsm fsm_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
fsm fsm_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
fsm fsm_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
fsm fsm_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
fsm fsm_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
fsm fsm_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
fsm fsm_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
xor_module xor_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
xor_module xor_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
fsm fsm_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
xor_module xor_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
xor_module xor_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
fsm fsm_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
fsm fsm_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
fsm fsm_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
xor_module xor_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
fsm fsm_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
xor_module xor_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
xor_module xor_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
fsm fsm_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
fsm fsm_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
xor_module xor_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
fsm fsm_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
xor_module xor_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
fsm fsm_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
fsm fsm_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
fsm fsm_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
fsm fsm_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
xor_module xor_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
fsm fsm_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
fsm fsm_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
fsm fsm_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
xor_module xor_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
fsm fsm_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
fsm fsm_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
xor_module xor_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
fsm fsm_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
fsm fsm_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
xor_module xor_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
fsm fsm_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
xor_module xor_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
fsm fsm_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
xor_module xor_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
fsm fsm_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
fsm fsm_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
xor_module xor_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
xor_module xor_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
xor_module xor_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
xor_module xor_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
fsm fsm_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
xor_module xor_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
fsm fsm_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
fsm fsm_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
fsm fsm_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
xor_module xor_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
fsm fsm_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
xor_module xor_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
xor_module xor_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
xor_module xor_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
xor_module xor_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
xor_module xor_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
fsm fsm_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
fsm fsm_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
fsm fsm_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
fsm fsm_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
xor_module xor_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
fsm fsm_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
fsm fsm_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
fsm fsm_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
fsm fsm_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
xor_module xor_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
fsm fsm_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
fsm fsm_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
fsm fsm_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
xor_module xor_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
fsm fsm_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
fsm fsm_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
fsm fsm_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
xor_module xor_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
xor_module xor_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
fsm fsm_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
fsm fsm_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
xor_module xor_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
xor_module xor_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
fsm fsm_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
fsm fsm_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
fsm fsm_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
fsm fsm_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
fsm fsm_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
fsm fsm_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
fsm fsm_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
fsm fsm_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
xor_module xor_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
xor_module xor_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
fsm fsm_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
fsm fsm_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
xor_module xor_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
fsm fsm_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
xor_module xor_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
fsm fsm_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
xor_module xor_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
fsm fsm_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
xor_module xor_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
xor_module xor_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
fsm fsm_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
fsm fsm_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
fsm fsm_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
fsm fsm_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
xor_module xor_module_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
xor_module xor_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
xor_module xor_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
xor_module xor_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
xor_module xor_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
fsm fsm_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
xor_module xor_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
xor_module xor_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
xor_module xor_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
fsm fsm_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
fsm fsm_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
fsm fsm_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
fsm fsm_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
xor_module xor_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
fsm fsm_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
xor_module xor_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
xor_module xor_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
fsm fsm_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
xor_module xor_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
fsm fsm_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
fsm fsm_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
fsm fsm_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
fsm fsm_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
xor_module xor_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
xor_module xor_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
fsm fsm_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
xor_module xor_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
fsm fsm_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
xor_module xor_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
xor_module xor_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
fsm fsm_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
fsm fsm_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
fsm fsm_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
xor_module xor_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
xor_module xor_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
xor_module xor_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
xor_module xor_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
xor_module xor_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
fsm fsm_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
xor_module xor_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
fsm fsm_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
fsm fsm_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
xor_module xor_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
fsm fsm_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
xor_module xor_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
fsm fsm_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
xor_module xor_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
fsm fsm_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
fsm fsm_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
fsm fsm_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
xor_module xor_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
xor_module xor_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
fsm fsm_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
fsm fsm_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
fsm fsm_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
fsm fsm_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
fsm fsm_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
xor_module xor_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
xor_module xor_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
fsm fsm_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
xor_module xor_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
xor_module xor_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
xor_module xor_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
xor_module xor_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
xor_module xor_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
xor_module xor_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
xor_module xor_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
fsm fsm_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
xor_module xor_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
fsm fsm_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
fsm fsm_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
fsm fsm_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
fsm fsm_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
fsm fsm_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
fsm fsm_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
fsm fsm_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
xor_module xor_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
xor_module xor_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
xor_module xor_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
fsm fsm_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
fsm fsm_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
fsm fsm_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
xor_module xor_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
xor_module xor_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
fsm fsm_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
xor_module xor_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
xor_module xor_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
xor_module xor_module_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
fsm fsm_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
fsm fsm_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
xor_module xor_module_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
fsm fsm_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
fsm fsm_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
xor_module xor_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
xor_module xor_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
xor_module xor_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
xor_module xor_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
xor_module xor_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
fsm fsm_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
fsm fsm_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
fsm fsm_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
fsm fsm_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
fsm fsm_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
fsm fsm_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
xor_module xor_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
fsm fsm_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
fsm fsm_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
xor_module xor_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
fsm fsm_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
fsm fsm_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
xor_module xor_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
fsm fsm_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
fsm fsm_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
xor_module xor_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
xor_module xor_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
xor_module xor_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
fsm fsm_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
fsm fsm_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
fsm fsm_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
xor_module xor_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
fsm fsm_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
xor_module xor_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
fsm fsm_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
fsm fsm_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
fsm fsm_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
fsm fsm_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
xor_module xor_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
xor_module xor_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
fsm fsm_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
fsm fsm_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
fsm fsm_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
xor_module xor_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
xor_module xor_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
fsm fsm_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
fsm fsm_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
fsm fsm_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
fsm fsm_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
fsm fsm_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
fsm fsm_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
fsm fsm_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
fsm fsm_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
fsm fsm_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
xor_module xor_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
xor_module xor_module_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
xor_module xor_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
xor_module xor_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
fsm fsm_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
xor_module xor_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
fsm fsm_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
fsm fsm_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
fsm fsm_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
xor_module xor_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
fsm fsm_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
xor_module xor_module_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
xor_module xor_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
xor_module xor_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
fsm fsm_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
fsm fsm_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
fsm fsm_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
fsm fsm_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
xor_module xor_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
fsm fsm_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
fsm fsm_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
xor_module xor_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
fsm fsm_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
xor_module xor_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
xor_module xor_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
fsm fsm_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
fsm fsm_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
fsm fsm_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
xor_module xor_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
xor_module xor_module_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
xor_module xor_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
fsm fsm_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
fsm fsm_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
fsm fsm_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [1157:0] <= intermediate_reg_1; 
outp[2119:1158] <= intermediate_reg_1[961:0] ; 
end 
endmodule 
 

module interface_4(input [331:0] inp, output reg [1775:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[331:0] <= inp ; 
outp[663:332] <= inp ; 
outp[995:664] <= inp ; 
outp[1327:996] <= inp ; 
outp[1659:1328] <= inp ; 
outp[1775:1660] <= inp[115:0] ; 
end 
endmodule 

module interface_5(input [1003:0] inp, output reg [1031:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[1003:0] <= inp ; 
outp[1031:1004] <= inp[27:0] ; 
end 
endmodule 

module interface_6(input [1003:0] inp, output reg [2519:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[1003:0] <= inp ; 
outp[2007:1004] <= inp ; 
outp[2519:2008] <= inp[511:0] ; 
end 
endmodule 

module interface_7(input [2007:0] inp, output reg [1133:0] outp, input clk, input reset);
reg [2007:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1003:0]intermediate_reg_1; 
 
xor_module xor_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
fsm fsm_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001])); 
fsm fsm_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
xor_module xor_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
fsm fsm_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
xor_module xor_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
fsm fsm_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
xor_module xor_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
fsm fsm_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
fsm fsm_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
fsm fsm_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
fsm fsm_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
fsm fsm_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
fsm fsm_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
xor_module xor_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
fsm fsm_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978])); 
fsm fsm_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
xor_module xor_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975])); 
fsm fsm_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974])); 
xor_module xor_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
xor_module xor_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
xor_module xor_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
fsm fsm_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
fsm fsm_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
xor_module xor_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
fsm fsm_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959])); 
xor_module xor_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
fsm fsm_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
fsm fsm_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
xor_module xor_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954])); 
fsm fsm_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
xor_module xor_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
fsm fsm_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950])); 
fsm fsm_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
fsm fsm_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948])); 
fsm fsm_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
xor_module xor_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
fsm fsm_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
fsm fsm_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
fsm fsm_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
fsm fsm_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
fsm fsm_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
fsm fsm_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
xor_module xor_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
fsm fsm_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
fsm fsm_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
fsm fsm_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
fsm fsm_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
fsm fsm_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
xor_module xor_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
xor_module xor_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
fsm fsm_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
fsm fsm_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
fsm fsm_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
fsm fsm_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
fsm fsm_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
fsm fsm_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
xor_module xor_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
fsm fsm_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906])); 
fsm fsm_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
fsm fsm_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
fsm fsm_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
fsm fsm_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
xor_module xor_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
fsm fsm_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
fsm fsm_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
fsm fsm_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
fsm fsm_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
xor_module xor_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884])); 
fsm fsm_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
xor_module xor_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
xor_module xor_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
fsm fsm_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
xor_module xor_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
xor_module xor_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
xor_module xor_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
fsm fsm_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
fsm fsm_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
xor_module xor_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
xor_module xor_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
xor_module xor_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
fsm fsm_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
xor_module xor_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
fsm fsm_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
xor_module xor_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
fsm fsm_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
fsm fsm_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
fsm fsm_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842])); 
xor_module xor_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
fsm fsm_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
xor_module xor_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
fsm fsm_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
xor_module xor_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
fsm fsm_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831])); 
fsm fsm_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829])); 
fsm fsm_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
fsm fsm_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
fsm fsm_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
fsm fsm_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823])); 
fsm fsm_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
fsm fsm_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
fsm fsm_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
xor_module xor_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
fsm fsm_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
xor_module xor_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
xor_module xor_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
fsm fsm_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
fsm fsm_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
fsm fsm_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
fsm fsm_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810])); 
xor_module xor_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
xor_module xor_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
fsm fsm_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
xor_module xor_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
xor_module xor_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
xor_module xor_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
xor_module xor_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
xor_module xor_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
fsm fsm_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
fsm fsm_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
fsm fsm_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
fsm fsm_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
fsm fsm_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
xor_module xor_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
xor_module xor_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
xor_module xor_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
xor_module xor_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
fsm fsm_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
xor_module xor_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
fsm fsm_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
fsm fsm_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
fsm fsm_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
fsm fsm_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
xor_module xor_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
fsm fsm_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
xor_module xor_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
xor_module xor_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
xor_module xor_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
fsm fsm_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
fsm fsm_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
xor_module xor_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
xor_module xor_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
xor_module xor_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
fsm fsm_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
xor_module xor_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
fsm fsm_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
xor_module xor_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
fsm fsm_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
xor_module xor_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
fsm fsm_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
xor_module xor_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
fsm fsm_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
fsm fsm_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
fsm fsm_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
xor_module xor_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
xor_module xor_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
fsm fsm_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
xor_module xor_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
xor_module xor_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
fsm fsm_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
fsm fsm_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
xor_module xor_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
xor_module xor_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
xor_module xor_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
fsm fsm_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
fsm fsm_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
xor_module xor_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
fsm fsm_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
xor_module xor_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
xor_module xor_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
fsm fsm_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
fsm fsm_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
fsm fsm_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
xor_module xor_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
xor_module xor_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
fsm fsm_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
fsm fsm_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
fsm fsm_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
fsm fsm_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
fsm fsm_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
fsm fsm_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
fsm fsm_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
fsm fsm_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
fsm fsm_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
fsm fsm_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
fsm fsm_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687])); 
xor_module xor_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
fsm fsm_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
fsm fsm_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
xor_module xor_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
xor_module xor_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
xor_module xor_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
fsm fsm_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
fsm fsm_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
fsm fsm_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
fsm fsm_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
fsm fsm_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
fsm fsm_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
xor_module xor_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
fsm fsm_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
fsm fsm_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
fsm fsm_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
fsm fsm_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
fsm fsm_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
fsm fsm_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
fsm fsm_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
fsm fsm_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
xor_module xor_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
xor_module xor_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
xor_module xor_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
fsm fsm_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
fsm fsm_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
fsm fsm_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
fsm fsm_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
fsm fsm_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
xor_module xor_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
xor_module xor_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
fsm fsm_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
fsm fsm_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
fsm fsm_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
xor_module xor_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
fsm fsm_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
fsm fsm_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
fsm fsm_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
xor_module xor_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
fsm fsm_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
fsm fsm_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
fsm fsm_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
xor_module xor_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
xor_module xor_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
fsm fsm_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
fsm fsm_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
fsm fsm_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
xor_module xor_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
fsm fsm_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
fsm fsm_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
fsm fsm_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
fsm fsm_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
fsm fsm_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
xor_module xor_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
xor_module xor_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
fsm fsm_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
fsm fsm_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
xor_module xor_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
fsm fsm_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
xor_module xor_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
xor_module xor_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
xor_module xor_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
fsm fsm_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
fsm fsm_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
fsm fsm_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
xor_module xor_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
xor_module xor_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
fsm fsm_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
xor_module xor_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
fsm fsm_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
fsm fsm_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
fsm fsm_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
fsm fsm_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
xor_module xor_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
fsm fsm_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
fsm fsm_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
fsm fsm_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
xor_module xor_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
fsm fsm_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
fsm fsm_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
fsm fsm_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
fsm fsm_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
fsm fsm_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
fsm fsm_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
xor_module xor_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
fsm fsm_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
xor_module xor_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
xor_module xor_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
fsm fsm_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
xor_module xor_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
fsm fsm_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
xor_module xor_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
xor_module xor_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
xor_module xor_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
xor_module xor_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
fsm fsm_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
fsm fsm_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
fsm fsm_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
fsm fsm_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
xor_module xor_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
xor_module xor_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
fsm fsm_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
xor_module xor_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
fsm fsm_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
fsm fsm_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
fsm fsm_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
xor_module xor_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
fsm fsm_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
xor_module xor_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
fsm fsm_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
fsm fsm_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
xor_module xor_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
fsm fsm_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
fsm fsm_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
xor_module xor_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
xor_module xor_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
xor_module xor_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
fsm fsm_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
xor_module xor_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
xor_module xor_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
fsm fsm_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
xor_module xor_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
xor_module xor_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
xor_module xor_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
fsm fsm_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
fsm fsm_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
fsm fsm_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
xor_module xor_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
fsm fsm_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
fsm fsm_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
xor_module xor_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
xor_module xor_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
xor_module xor_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
fsm fsm_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
fsm fsm_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
fsm fsm_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
fsm fsm_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
fsm fsm_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
fsm fsm_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
xor_module xor_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
xor_module xor_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
fsm fsm_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
fsm fsm_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
xor_module xor_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
xor_module xor_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
fsm fsm_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
xor_module xor_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
fsm fsm_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
xor_module xor_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
xor_module xor_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
xor_module xor_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
fsm fsm_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
fsm fsm_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
fsm fsm_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
fsm fsm_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
xor_module xor_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
xor_module xor_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
fsm fsm_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
fsm fsm_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
fsm fsm_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
fsm fsm_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
xor_module xor_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
xor_module xor_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
fsm fsm_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
xor_module xor_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
fsm fsm_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
fsm fsm_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
xor_module xor_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
fsm fsm_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
fsm fsm_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
fsm fsm_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
fsm fsm_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
fsm fsm_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
xor_module xor_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
fsm fsm_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
xor_module xor_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
xor_module xor_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
xor_module xor_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
fsm fsm_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
xor_module xor_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
fsm fsm_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
xor_module xor_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
fsm fsm_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
xor_module xor_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
fsm fsm_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
fsm fsm_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
fsm fsm_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
fsm fsm_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
xor_module xor_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
xor_module xor_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
xor_module xor_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
fsm fsm_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
xor_module xor_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
xor_module xor_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
xor_module xor_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
xor_module xor_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
xor_module xor_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
fsm fsm_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
xor_module xor_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
xor_module xor_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
fsm fsm_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
fsm fsm_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
fsm fsm_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
xor_module xor_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
fsm fsm_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
xor_module xor_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
fsm fsm_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
fsm fsm_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
xor_module xor_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
xor_module xor_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
fsm fsm_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
xor_module xor_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
fsm fsm_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
fsm fsm_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
xor_module xor_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
fsm fsm_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
fsm fsm_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
fsm fsm_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
xor_module xor_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
fsm fsm_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
fsm fsm_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
xor_module xor_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
xor_module xor_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
xor_module xor_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
xor_module xor_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
fsm fsm_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
xor_module xor_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
xor_module xor_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
fsm fsm_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
fsm fsm_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
xor_module xor_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
fsm fsm_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
xor_module xor_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
xor_module xor_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
xor_module xor_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
xor_module xor_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
xor_module xor_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
xor_module xor_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
xor_module xor_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
fsm fsm_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
xor_module xor_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
xor_module xor_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
xor_module xor_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
fsm fsm_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
xor_module xor_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
xor_module xor_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
xor_module xor_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
fsm fsm_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
fsm fsm_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
xor_module xor_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
fsm fsm_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
xor_module xor_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
xor_module xor_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
xor_module xor_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
fsm fsm_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
fsm fsm_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
fsm fsm_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
fsm fsm_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
xor_module xor_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
fsm fsm_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
fsm fsm_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
xor_module xor_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
xor_module xor_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
fsm fsm_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
xor_module xor_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
xor_module xor_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
fsm fsm_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
xor_module xor_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
xor_module xor_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
fsm fsm_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
fsm fsm_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
fsm fsm_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
xor_module xor_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
xor_module xor_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
fsm fsm_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
fsm fsm_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
fsm fsm_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
fsm fsm_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
xor_module xor_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
xor_module xor_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
fsm fsm_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
xor_module xor_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
fsm fsm_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
fsm fsm_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
fsm fsm_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
xor_module xor_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
fsm fsm_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
fsm fsm_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
xor_module xor_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
fsm fsm_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
fsm fsm_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
xor_module xor_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
xor_module xor_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
xor_module xor_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
xor_module xor_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
fsm fsm_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
fsm fsm_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
xor_module xor_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
fsm fsm_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
xor_module xor_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
xor_module xor_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
xor_module xor_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
fsm fsm_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
fsm fsm_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
fsm fsm_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
xor_module xor_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
xor_module xor_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
fsm fsm_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
fsm fsm_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
xor_module xor_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
xor_module xor_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
xor_module xor_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
fsm fsm_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
xor_module xor_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
fsm fsm_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
fsm fsm_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
xor_module xor_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
xor_module xor_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
xor_module xor_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
fsm fsm_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
xor_module xor_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
xor_module xor_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
fsm fsm_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
xor_module xor_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
fsm fsm_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
xor_module xor_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
fsm fsm_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
xor_module xor_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
fsm fsm_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
fsm fsm_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
fsm fsm_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
xor_module xor_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
xor_module xor_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
fsm fsm_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
fsm fsm_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
fsm fsm_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
fsm fsm_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
xor_module xor_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
xor_module xor_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
xor_module xor_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
xor_module xor_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
fsm fsm_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
xor_module xor_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
fsm fsm_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
xor_module xor_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
fsm fsm_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
fsm fsm_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
fsm fsm_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
xor_module xor_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
xor_module xor_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
xor_module xor_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
xor_module xor_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
fsm fsm_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
fsm fsm_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
fsm fsm_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
fsm fsm_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
fsm fsm_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
xor_module xor_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
xor_module xor_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
xor_module xor_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
xor_module xor_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
fsm fsm_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
fsm fsm_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
fsm fsm_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
xor_module xor_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
fsm fsm_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
fsm fsm_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
fsm fsm_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
xor_module xor_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
xor_module xor_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
fsm fsm_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
xor_module xor_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
fsm fsm_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
fsm fsm_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
xor_module xor_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
fsm fsm_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
xor_module xor_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
fsm fsm_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
fsm fsm_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
xor_module xor_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
xor_module xor_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
xor_module xor_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
fsm fsm_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
xor_module xor_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
xor_module xor_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
xor_module xor_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
xor_module xor_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
fsm fsm_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
xor_module xor_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
xor_module xor_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
xor_module xor_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
fsm fsm_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
xor_module xor_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
xor_module xor_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
xor_module xor_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
xor_module xor_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
xor_module xor_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
xor_module xor_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
fsm fsm_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
fsm fsm_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
fsm fsm_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
fsm fsm_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
xor_module xor_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
xor_module xor_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
fsm fsm_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
xor_module xor_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
fsm fsm_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
xor_module xor_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
xor_module xor_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
xor_module xor_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
fsm fsm_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
xor_module xor_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
xor_module xor_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
xor_module xor_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
fsm fsm_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
xor_module xor_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
fsm fsm_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
fsm fsm_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
fsm fsm_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
xor_module xor_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
fsm fsm_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
fsm fsm_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
xor_module xor_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
fsm fsm_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
fsm fsm_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
xor_module xor_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
xor_module xor_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
fsm fsm_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
fsm fsm_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
fsm fsm_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
xor_module xor_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
fsm fsm_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
fsm fsm_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
fsm fsm_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
xor_module xor_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
xor_module xor_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
fsm fsm_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
xor_module xor_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
xor_module xor_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
xor_module xor_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
fsm fsm_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
fsm fsm_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
xor_module xor_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
xor_module xor_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
fsm fsm_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
fsm fsm_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
xor_module xor_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
xor_module xor_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
xor_module xor_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
fsm fsm_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
fsm fsm_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
fsm fsm_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
fsm fsm_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
xor_module xor_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
xor_module xor_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
xor_module xor_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
xor_module xor_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
xor_module xor_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
fsm fsm_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
fsm fsm_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
fsm fsm_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
fsm fsm_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
xor_module xor_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
xor_module xor_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
xor_module xor_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
fsm fsm_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
xor_module xor_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
xor_module xor_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
xor_module xor_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
xor_module xor_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
fsm fsm_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
xor_module xor_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
fsm fsm_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
fsm fsm_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
fsm fsm_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
fsm fsm_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
xor_module xor_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
xor_module xor_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
fsm fsm_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
xor_module xor_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
xor_module xor_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
fsm fsm_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
fsm fsm_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
fsm fsm_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
xor_module xor_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
fsm fsm_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
xor_module xor_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
xor_module xor_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
fsm fsm_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
fsm fsm_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
xor_module xor_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
fsm fsm_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
xor_module xor_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
fsm fsm_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
fsm fsm_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
fsm fsm_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
xor_module xor_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
fsm fsm_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [1003:0] <= intermediate_reg_1; 
outp[1133:1004] <= intermediate_reg_1[129:0] ; 
end 
endmodule 
 

module interface_8(input [2007:0] inp, output reg [1117:0] outp, input clk, input reset);
reg [2007:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1003:0]intermediate_reg_1; 
 
fsm fsm_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
fsm fsm_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001])); 
fsm fsm_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
xor_module xor_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
xor_module xor_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
fsm fsm_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991])); 
fsm fsm_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
fsm fsm_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
xor_module xor_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
fsm fsm_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
xor_module xor_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
fsm fsm_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
fsm fsm_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
fsm fsm_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
xor_module xor_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
fsm fsm_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
fsm fsm_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
fsm fsm_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
xor_module xor_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974])); 
fsm fsm_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
xor_module xor_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
fsm fsm_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971])); 
fsm fsm_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
fsm fsm_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
fsm fsm_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
fsm fsm_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962])); 
fsm fsm_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959])); 
fsm fsm_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
fsm fsm_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
fsm fsm_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954])); 
fsm fsm_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
fsm fsm_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
xor_module xor_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
xor_module xor_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950])); 
fsm fsm_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
fsm fsm_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
fsm fsm_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
xor_module xor_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
fsm fsm_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
fsm fsm_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
fsm fsm_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
fsm fsm_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
xor_module xor_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
xor_module xor_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
xor_module xor_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
xor_module xor_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
fsm fsm_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
xor_module xor_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
fsm fsm_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
fsm fsm_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
fsm fsm_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
fsm fsm_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
fsm fsm_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
fsm fsm_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
fsm fsm_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
fsm fsm_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
xor_module xor_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
xor_module xor_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
xor_module xor_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
xor_module xor_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
fsm fsm_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
xor_module xor_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
fsm fsm_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
fsm fsm_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
fsm fsm_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
fsm fsm_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
fsm fsm_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
xor_module xor_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884])); 
xor_module xor_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
fsm fsm_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
xor_module xor_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
xor_module xor_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
fsm fsm_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
fsm fsm_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
fsm fsm_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
fsm fsm_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
fsm fsm_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
fsm fsm_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
fsm fsm_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
xor_module xor_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862])); 
fsm fsm_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
fsm fsm_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
fsm fsm_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
fsm fsm_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
xor_module xor_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
xor_module xor_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
fsm fsm_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
fsm fsm_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
fsm fsm_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
fsm fsm_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842])); 
xor_module xor_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
fsm fsm_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
fsm fsm_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
fsm fsm_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
fsm fsm_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
fsm fsm_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831])); 
fsm fsm_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829])); 
fsm fsm_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
fsm fsm_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823])); 
xor_module xor_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
fsm fsm_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
xor_module xor_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
fsm fsm_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
xor_module xor_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
fsm fsm_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
fsm fsm_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
fsm fsm_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
fsm fsm_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
fsm fsm_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810])); 
fsm fsm_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
xor_module xor_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
fsm fsm_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
xor_module xor_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
fsm fsm_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
fsm fsm_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
fsm fsm_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
xor_module xor_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
xor_module xor_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
fsm fsm_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
xor_module xor_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
fsm fsm_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
fsm fsm_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
fsm fsm_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
xor_module xor_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
fsm fsm_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
xor_module xor_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
fsm fsm_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
fsm fsm_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
fsm fsm_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
fsm fsm_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
fsm fsm_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
fsm fsm_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
xor_module xor_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
xor_module xor_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
fsm fsm_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
fsm fsm_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
fsm fsm_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
fsm fsm_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
xor_module xor_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
xor_module xor_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
fsm fsm_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
fsm fsm_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
fsm fsm_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
fsm fsm_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
xor_module xor_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
fsm fsm_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
fsm fsm_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
xor_module xor_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
xor_module xor_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
fsm fsm_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
xor_module xor_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
fsm fsm_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
xor_module xor_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
fsm fsm_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
fsm fsm_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
fsm fsm_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
fsm fsm_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
xor_module xor_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
xor_module xor_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
fsm fsm_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
fsm fsm_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
xor_module xor_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
xor_module xor_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
fsm fsm_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
xor_module xor_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
fsm fsm_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
xor_module xor_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
fsm fsm_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
fsm fsm_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
xor_module xor_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
fsm fsm_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
fsm fsm_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
xor_module xor_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
fsm fsm_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
fsm fsm_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
fsm fsm_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
fsm fsm_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
fsm fsm_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
fsm fsm_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
fsm fsm_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
fsm fsm_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
fsm fsm_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687])); 
fsm fsm_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
fsm fsm_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
fsm fsm_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
xor_module xor_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
fsm fsm_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
xor_module xor_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
fsm fsm_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
xor_module xor_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
fsm fsm_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
fsm fsm_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
xor_module xor_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
fsm fsm_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
fsm fsm_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
fsm fsm_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
fsm fsm_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
xor_module xor_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
fsm fsm_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
fsm fsm_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
fsm fsm_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
fsm fsm_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
fsm fsm_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
fsm fsm_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
fsm fsm_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
fsm fsm_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
xor_module xor_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
fsm fsm_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
fsm fsm_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
xor_module xor_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
fsm fsm_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
fsm fsm_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
xor_module xor_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
fsm fsm_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
fsm fsm_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
fsm fsm_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
fsm fsm_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
fsm fsm_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
xor_module xor_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
xor_module xor_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
xor_module xor_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
fsm fsm_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
xor_module xor_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
fsm fsm_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
fsm fsm_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
xor_module xor_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
xor_module xor_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
fsm fsm_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
xor_module xor_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
fsm fsm_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
xor_module xor_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
fsm fsm_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
fsm fsm_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
xor_module xor_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
xor_module xor_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
xor_module xor_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
fsm fsm_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
xor_module xor_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
fsm fsm_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
fsm fsm_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
fsm fsm_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
fsm fsm_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
xor_module xor_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
fsm fsm_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
fsm fsm_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
xor_module xor_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
fsm fsm_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
fsm fsm_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
xor_module xor_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
fsm fsm_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
fsm fsm_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
xor_module xor_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
xor_module xor_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
fsm fsm_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
fsm fsm_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
fsm fsm_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
fsm fsm_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
fsm fsm_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
fsm fsm_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
xor_module xor_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
xor_module xor_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
xor_module xor_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
fsm fsm_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
xor_module xor_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
xor_module xor_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
xor_module xor_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
xor_module xor_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
xor_module xor_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
xor_module xor_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
xor_module xor_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
fsm fsm_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
fsm fsm_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
fsm fsm_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
xor_module xor_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
xor_module xor_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
fsm fsm_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
fsm fsm_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
xor_module xor_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
xor_module xor_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
fsm fsm_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
fsm fsm_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
xor_module xor_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
fsm fsm_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
fsm fsm_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
fsm fsm_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
fsm fsm_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
fsm fsm_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
xor_module xor_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
xor_module xor_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
fsm fsm_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
fsm fsm_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
xor_module xor_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
xor_module xor_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
fsm fsm_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
fsm fsm_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
xor_module xor_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
xor_module xor_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
fsm fsm_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
xor_module xor_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
xor_module xor_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
fsm fsm_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
fsm fsm_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
fsm fsm_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
xor_module xor_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
xor_module xor_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
xor_module xor_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
fsm fsm_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
xor_module xor_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
fsm fsm_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
fsm fsm_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
xor_module xor_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
fsm fsm_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
fsm fsm_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
xor_module xor_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
fsm fsm_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
fsm fsm_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
xor_module xor_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
fsm fsm_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
fsm fsm_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
xor_module xor_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
xor_module xor_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
xor_module xor_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
fsm fsm_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
xor_module xor_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
fsm fsm_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
fsm fsm_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
fsm fsm_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
xor_module xor_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
xor_module xor_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
fsm fsm_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
fsm fsm_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
fsm fsm_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
fsm fsm_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
fsm fsm_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
fsm fsm_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
fsm fsm_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
fsm fsm_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
fsm fsm_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
fsm fsm_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
fsm fsm_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
fsm fsm_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
fsm fsm_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
xor_module xor_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
xor_module xor_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
fsm fsm_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
xor_module xor_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
fsm fsm_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
xor_module xor_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
fsm fsm_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
xor_module xor_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
fsm fsm_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
fsm fsm_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
fsm fsm_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
fsm fsm_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
xor_module xor_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
xor_module xor_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
xor_module xor_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
xor_module xor_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
xor_module xor_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
fsm fsm_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
fsm fsm_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
fsm fsm_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
xor_module xor_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
fsm fsm_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
fsm fsm_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
fsm fsm_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
xor_module xor_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
xor_module xor_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
fsm fsm_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
xor_module xor_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
fsm fsm_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
xor_module xor_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
xor_module xor_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
fsm fsm_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
xor_module xor_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
xor_module xor_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
fsm fsm_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
xor_module xor_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
xor_module xor_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
xor_module xor_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
fsm fsm_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
xor_module xor_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
xor_module xor_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
fsm fsm_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
xor_module xor_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
xor_module xor_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
xor_module xor_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
xor_module xor_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
fsm fsm_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
fsm fsm_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
fsm fsm_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
fsm fsm_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
fsm fsm_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
fsm fsm_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
xor_module xor_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
xor_module xor_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
xor_module xor_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
xor_module xor_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
fsm fsm_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
fsm fsm_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
fsm fsm_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
fsm fsm_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
fsm fsm_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
fsm fsm_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
fsm fsm_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
fsm fsm_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
fsm fsm_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
fsm fsm_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
fsm fsm_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
fsm fsm_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
xor_module xor_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
fsm fsm_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
xor_module xor_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
fsm fsm_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
xor_module xor_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
xor_module xor_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
fsm fsm_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
fsm fsm_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
fsm fsm_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
fsm fsm_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
fsm fsm_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
xor_module xor_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
fsm fsm_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
xor_module xor_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
fsm fsm_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
xor_module xor_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
fsm fsm_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
fsm fsm_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
fsm fsm_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
xor_module xor_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
fsm fsm_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
xor_module xor_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
xor_module xor_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
xor_module xor_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
fsm fsm_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
xor_module xor_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
fsm fsm_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
fsm fsm_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
fsm fsm_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
fsm fsm_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
fsm fsm_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
xor_module xor_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
fsm fsm_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
fsm fsm_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
fsm fsm_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
xor_module xor_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
xor_module xor_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
fsm fsm_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
xor_module xor_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
fsm fsm_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
xor_module xor_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
fsm fsm_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
fsm fsm_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
fsm fsm_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
fsm fsm_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
fsm fsm_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
fsm fsm_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
xor_module xor_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
fsm fsm_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
xor_module xor_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
fsm fsm_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
xor_module xor_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
fsm fsm_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
xor_module xor_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
fsm fsm_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
xor_module xor_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
xor_module xor_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
fsm fsm_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
xor_module xor_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
fsm fsm_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
fsm fsm_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
fsm fsm_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
xor_module xor_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
xor_module xor_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
fsm fsm_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
xor_module xor_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
xor_module xor_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
xor_module xor_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
fsm fsm_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
xor_module xor_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
xor_module xor_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
fsm fsm_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
fsm fsm_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
fsm fsm_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
xor_module xor_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
xor_module xor_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
fsm fsm_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
xor_module xor_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
xor_module xor_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
xor_module xor_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
xor_module xor_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
xor_module xor_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
xor_module xor_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
xor_module xor_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
xor_module xor_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
fsm fsm_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
fsm fsm_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
xor_module xor_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
fsm fsm_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
fsm fsm_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
fsm fsm_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
fsm fsm_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
xor_module xor_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
fsm fsm_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
xor_module xor_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
fsm fsm_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
xor_module xor_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
fsm fsm_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
fsm fsm_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
xor_module xor_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
xor_module xor_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
fsm fsm_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
xor_module xor_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
xor_module xor_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
xor_module xor_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
fsm fsm_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
xor_module xor_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
fsm fsm_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
xor_module xor_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
xor_module xor_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
xor_module xor_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
fsm fsm_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
fsm fsm_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
xor_module xor_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
fsm fsm_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
xor_module xor_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
fsm fsm_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
xor_module xor_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
fsm fsm_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
xor_module xor_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
fsm fsm_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
xor_module xor_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
xor_module xor_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
xor_module xor_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
fsm fsm_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
fsm fsm_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
fsm fsm_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
fsm fsm_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
fsm fsm_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
fsm fsm_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
xor_module xor_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
xor_module xor_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
xor_module xor_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
fsm fsm_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
xor_module xor_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
xor_module xor_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
xor_module xor_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
xor_module xor_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
fsm fsm_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
xor_module xor_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
fsm fsm_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
xor_module xor_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
xor_module xor_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
xor_module xor_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
fsm fsm_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
xor_module xor_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
fsm fsm_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
fsm fsm_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
fsm fsm_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
fsm fsm_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
xor_module xor_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
fsm fsm_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
xor_module xor_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
fsm fsm_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
fsm fsm_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
xor_module xor_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
xor_module xor_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
fsm fsm_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
xor_module xor_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
xor_module xor_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
xor_module xor_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
xor_module xor_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
xor_module xor_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
xor_module xor_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
fsm fsm_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
fsm fsm_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
xor_module xor_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
xor_module xor_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
fsm fsm_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
fsm fsm_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
fsm fsm_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
fsm fsm_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
fsm fsm_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
fsm fsm_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
xor_module xor_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
xor_module xor_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
xor_module xor_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
fsm fsm_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
fsm fsm_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
fsm fsm_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
fsm fsm_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
xor_module xor_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
xor_module xor_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
xor_module xor_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
fsm fsm_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
fsm fsm_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
fsm fsm_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
xor_module xor_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
fsm fsm_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
fsm fsm_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
xor_module xor_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
xor_module xor_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
xor_module xor_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
fsm fsm_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
fsm fsm_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
xor_module xor_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
xor_module xor_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
fsm fsm_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
xor_module xor_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
xor_module xor_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
fsm fsm_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
fsm fsm_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
fsm fsm_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
xor_module xor_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
fsm fsm_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
fsm fsm_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
xor_module xor_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
fsm fsm_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
xor_module xor_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
xor_module xor_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
xor_module xor_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
xor_module xor_module_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
xor_module xor_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
fsm fsm_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
fsm fsm_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
xor_module xor_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
fsm fsm_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
fsm fsm_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
fsm fsm_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
xor_module xor_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
fsm fsm_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
xor_module xor_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
fsm fsm_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
fsm fsm_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
fsm fsm_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
xor_module xor_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
fsm fsm_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
fsm fsm_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
fsm fsm_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
xor_module xor_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
fsm fsm_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
fsm fsm_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
xor_module xor_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
fsm fsm_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
xor_module xor_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
xor_module xor_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
xor_module xor_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
fsm fsm_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
fsm fsm_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
xor_module xor_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
fsm fsm_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
fsm fsm_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
fsm fsm_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
fsm fsm_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
xor_module xor_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
fsm fsm_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
xor_module xor_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
fsm fsm_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
fsm fsm_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
xor_module xor_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
fsm fsm_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [1003:0] <= intermediate_reg_1; 
outp[1117:1004] <= intermediate_reg_1[113:0] ; 
end 
endmodule 
 

module interface_9(input [1007:0] inp, output reg [3551:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[1007:0] <= inp ; 
outp[2015:1008] <= inp ; 
outp[3023:2016] <= inp ; 
outp[3551:3024] <= inp[527:0] ; 
end 
endmodule 

module interface_10(input [2479:0] inp, output reg [1059:0] outp, input clk, input reset);
reg [2479:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1239:0]intermediate_reg_1; 
 
xor_module xor_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239])); 
xor_module xor_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236])); 
fsm fsm_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229])); 
xor_module xor_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227])); 
fsm fsm_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
fsm fsm_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225])); 
fsm fsm_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222])); 
fsm fsm_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
fsm fsm_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219])); 
fsm fsm_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218])); 
fsm fsm_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217])); 
fsm fsm_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215])); 
fsm fsm_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213])); 
fsm fsm_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212])); 
fsm fsm_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211])); 
fsm fsm_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210])); 
fsm fsm_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209])); 
fsm fsm_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208])); 
fsm fsm_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206])); 
fsm fsm_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204])); 
xor_module xor_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203])); 
fsm fsm_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202])); 
fsm fsm_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201])); 
fsm fsm_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197])); 
fsm fsm_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195])); 
fsm fsm_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191])); 
fsm fsm_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190])); 
fsm fsm_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189])); 
fsm fsm_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188])); 
fsm fsm_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187])); 
xor_module xor_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186])); 
xor_module xor_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183])); 
fsm fsm_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181])); 
fsm fsm_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178])); 
xor_module xor_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177])); 
fsm fsm_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174])); 
xor_module xor_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173])); 
fsm fsm_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172])); 
xor_module xor_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169])); 
xor_module xor_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168])); 
fsm fsm_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167])); 
xor_module xor_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166])); 
xor_module xor_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165])); 
fsm fsm_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163])); 
fsm fsm_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162])); 
fsm fsm_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161])); 
xor_module xor_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158])); 
fsm fsm_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156])); 
fsm fsm_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154])); 
fsm fsm_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152])); 
fsm fsm_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
fsm fsm_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146])); 
fsm fsm_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145])); 
fsm fsm_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143])); 
fsm fsm_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137])); 
fsm fsm_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136])); 
xor_module xor_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135])); 
xor_module xor_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134])); 
fsm fsm_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133])); 
fsm fsm_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129])); 
xor_module xor_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126])); 
xor_module xor_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
xor_module xor_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
fsm fsm_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120])); 
fsm fsm_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
fsm fsm_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118])); 
fsm fsm_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117])); 
fsm fsm_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114])); 
xor_module xor_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113])); 
xor_module xor_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112])); 
xor_module xor_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110])); 
xor_module xor_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
fsm fsm_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107])); 
fsm fsm_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106])); 
fsm fsm_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
xor_module xor_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
fsm fsm_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
fsm fsm_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102])); 
xor_module xor_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100])); 
fsm fsm_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099])); 
fsm fsm_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098])); 
fsm fsm_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096])); 
xor_module xor_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095])); 
fsm fsm_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094])); 
fsm fsm_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
fsm fsm_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
xor_module xor_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
xor_module xor_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
xor_module xor_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086])); 
fsm fsm_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085])); 
fsm fsm_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082])); 
fsm fsm_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
fsm fsm_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077])); 
xor_module xor_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
fsm fsm_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072])); 
fsm fsm_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
fsm fsm_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065])); 
xor_module xor_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061])); 
fsm fsm_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059])); 
fsm fsm_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057])); 
xor_module xor_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056])); 
xor_module xor_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055])); 
fsm fsm_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054])); 
fsm fsm_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053])); 
fsm fsm_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051])); 
fsm fsm_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050])); 
xor_module xor_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
xor_module xor_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046])); 
fsm fsm_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045])); 
fsm fsm_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
xor_module xor_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
xor_module xor_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041])); 
xor_module xor_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036])); 
fsm fsm_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034])); 
fsm fsm_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032])); 
fsm fsm_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
xor_module xor_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030])); 
xor_module xor_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029])); 
fsm fsm_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
fsm fsm_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027])); 
fsm fsm_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026])); 
xor_module xor_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
xor_module xor_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
fsm fsm_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
xor_module xor_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018])); 
xor_module xor_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017])); 
fsm fsm_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012])); 
fsm fsm_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011])); 
xor_module xor_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010])); 
xor_module xor_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
fsm fsm_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006])); 
fsm fsm_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
xor_module xor_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
xor_module xor_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
fsm fsm_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001])); 
fsm fsm_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
fsm fsm_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
fsm fsm_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
xor_module xor_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
xor_module xor_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991])); 
fsm fsm_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
fsm fsm_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
fsm fsm_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
fsm fsm_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
fsm fsm_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
xor_module xor_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
xor_module xor_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
fsm fsm_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
xor_module xor_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978])); 
xor_module xor_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
fsm fsm_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
fsm fsm_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975])); 
xor_module xor_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974])); 
xor_module xor_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970])); 
fsm fsm_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
xor_module xor_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
xor_module xor_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
fsm fsm_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
fsm fsm_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
xor_module xor_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959])); 
xor_module xor_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
fsm fsm_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
fsm fsm_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
xor_module xor_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
xor_module xor_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954])); 
fsm fsm_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
fsm fsm_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
fsm fsm_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948])); 
fsm fsm_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
xor_module xor_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
xor_module xor_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
fsm fsm_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
fsm fsm_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
fsm fsm_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
fsm fsm_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
fsm fsm_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
fsm fsm_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
xor_module xor_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
fsm fsm_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
fsm fsm_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
xor_module xor_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
fsm fsm_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
fsm fsm_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
xor_module xor_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
fsm fsm_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
fsm fsm_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
fsm fsm_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
fsm fsm_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
xor_module xor_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
fsm fsm_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
xor_module xor_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
fsm fsm_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
fsm fsm_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
fsm fsm_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
fsm fsm_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
fsm fsm_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
fsm fsm_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906])); 
fsm fsm_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
fsm fsm_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
fsm fsm_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
fsm fsm_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
fsm fsm_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
fsm fsm_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
fsm fsm_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
fsm fsm_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
fsm fsm_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
xor_module xor_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
xor_module xor_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
xor_module xor_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
fsm fsm_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
xor_module xor_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879])); 
fsm fsm_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
fsm fsm_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
fsm fsm_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
xor_module xor_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
fsm fsm_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
xor_module xor_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
xor_module xor_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
xor_module xor_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862])); 
fsm fsm_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
xor_module xor_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
xor_module xor_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
fsm fsm_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
fsm fsm_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
fsm fsm_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
xor_module xor_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
fsm fsm_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
fsm fsm_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
fsm fsm_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
fsm fsm_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
xor_module xor_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
fsm fsm_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
xor_module xor_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
fsm fsm_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
fsm fsm_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
fsm fsm_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
xor_module xor_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
fsm fsm_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831])); 
xor_module xor_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
fsm fsm_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
xor_module xor_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
xor_module xor_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
fsm fsm_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
fsm fsm_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
fsm fsm_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
fsm fsm_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
fsm fsm_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
xor_module xor_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
fsm fsm_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
xor_module xor_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
xor_module xor_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810])); 
fsm fsm_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
fsm fsm_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
xor_module xor_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
fsm fsm_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
xor_module xor_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
xor_module xor_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
xor_module xor_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
xor_module xor_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
fsm fsm_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
fsm fsm_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
fsm fsm_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
fsm fsm_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
xor_module xor_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
fsm fsm_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
fsm fsm_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
xor_module xor_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
fsm fsm_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
fsm fsm_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
fsm fsm_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
xor_module xor_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
fsm fsm_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
fsm fsm_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
xor_module xor_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
fsm fsm_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
fsm fsm_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
fsm fsm_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
xor_module xor_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
fsm fsm_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
xor_module xor_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
xor_module xor_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
xor_module xor_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
xor_module xor_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
xor_module xor_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
xor_module xor_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
xor_module xor_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
fsm fsm_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
fsm fsm_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
fsm fsm_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
fsm fsm_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
fsm fsm_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
fsm fsm_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
fsm fsm_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
fsm fsm_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
xor_module xor_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
fsm fsm_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
fsm fsm_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
fsm fsm_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
fsm fsm_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
fsm fsm_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
xor_module xor_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
xor_module xor_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
fsm fsm_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
fsm fsm_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
fsm fsm_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
fsm fsm_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
fsm fsm_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
xor_module xor_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
xor_module xor_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
xor_module xor_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
xor_module xor_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
xor_module xor_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
xor_module xor_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
xor_module xor_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
fsm fsm_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
fsm fsm_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
fsm fsm_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
xor_module xor_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
xor_module xor_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
fsm fsm_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
fsm fsm_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
xor_module xor_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
fsm fsm_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
fsm fsm_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
fsm fsm_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
xor_module xor_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
fsm fsm_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
xor_module xor_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
xor_module xor_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
fsm fsm_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
fsm fsm_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
fsm fsm_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
fsm fsm_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
fsm fsm_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687])); 
xor_module xor_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
fsm fsm_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
xor_module xor_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
fsm fsm_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
fsm fsm_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
xor_module xor_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
fsm fsm_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
xor_module xor_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
xor_module xor_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
xor_module xor_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
fsm fsm_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
xor_module xor_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
fsm fsm_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
xor_module xor_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
fsm fsm_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
fsm fsm_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
xor_module xor_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
fsm fsm_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
fsm fsm_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
fsm fsm_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
xor_module xor_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
xor_module xor_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
fsm fsm_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
fsm fsm_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
fsm fsm_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
xor_module xor_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642])); 
xor_module xor_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
xor_module xor_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640])); 
fsm fsm_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
fsm fsm_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
fsm fsm_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
fsm fsm_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
fsm fsm_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
fsm fsm_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
fsm fsm_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
fsm fsm_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
fsm fsm_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
fsm fsm_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
fsm fsm_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
fsm fsm_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
xor_module xor_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
xor_module xor_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
xor_module xor_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
xor_module xor_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
fsm fsm_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
xor_module xor_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
xor_module xor_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
xor_module xor_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
xor_module xor_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
xor_module xor_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
fsm fsm_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
xor_module xor_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
xor_module xor_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
fsm fsm_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
fsm fsm_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
xor_module xor_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
xor_module xor_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
fsm fsm_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
fsm fsm_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
fsm fsm_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
xor_module xor_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
fsm fsm_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
fsm fsm_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
fsm fsm_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
xor_module xor_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
fsm fsm_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
fsm fsm_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
fsm fsm_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
xor_module xor_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
xor_module xor_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
fsm fsm_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
fsm fsm_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
xor_module xor_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
fsm fsm_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
xor_module xor_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
fsm fsm_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
fsm fsm_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
xor_module xor_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
xor_module xor_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
fsm fsm_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
fsm fsm_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
xor_module xor_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
xor_module xor_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
xor_module xor_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
xor_module xor_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
fsm fsm_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
xor_module xor_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
xor_module xor_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
xor_module xor_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
xor_module xor_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
fsm fsm_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
xor_module xor_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
fsm fsm_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
xor_module xor_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
fsm fsm_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
fsm fsm_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
xor_module xor_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
fsm fsm_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
fsm fsm_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
fsm fsm_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
xor_module xor_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
xor_module xor_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
xor_module xor_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
xor_module xor_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
fsm fsm_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
fsm fsm_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
xor_module xor_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
xor_module xor_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
xor_module xor_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
fsm fsm_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
fsm fsm_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
fsm fsm_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
xor_module xor_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
fsm fsm_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
xor_module xor_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
fsm fsm_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
fsm fsm_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
xor_module xor_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
fsm fsm_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
xor_module xor_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
xor_module xor_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
fsm fsm_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
xor_module xor_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
xor_module xor_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
fsm fsm_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
fsm fsm_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
fsm fsm_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
xor_module xor_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
fsm fsm_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
fsm fsm_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
fsm fsm_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
fsm fsm_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
xor_module xor_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
fsm fsm_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
xor_module xor_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
xor_module xor_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
xor_module xor_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
xor_module xor_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
xor_module xor_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
xor_module xor_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
fsm fsm_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
fsm fsm_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
fsm fsm_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
fsm fsm_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
fsm fsm_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
xor_module xor_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
xor_module xor_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
fsm fsm_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
xor_module xor_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
fsm fsm_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
fsm fsm_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
xor_module xor_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
fsm fsm_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
xor_module xor_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
fsm fsm_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
xor_module xor_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
fsm fsm_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
xor_module xor_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
fsm fsm_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
xor_module xor_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
fsm fsm_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
xor_module xor_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
fsm fsm_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
xor_module xor_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
fsm fsm_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
fsm fsm_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
xor_module xor_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
fsm fsm_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
fsm fsm_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
xor_module xor_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
fsm fsm_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
xor_module xor_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
xor_module xor_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
xor_module xor_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
fsm fsm_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
fsm fsm_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
fsm fsm_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
fsm fsm_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
xor_module xor_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
xor_module xor_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
xor_module xor_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
xor_module xor_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
xor_module xor_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
fsm fsm_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
fsm fsm_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
xor_module xor_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
xor_module xor_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
fsm fsm_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
fsm fsm_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
fsm fsm_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
xor_module xor_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
fsm fsm_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
xor_module xor_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
fsm fsm_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
xor_module xor_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
xor_module xor_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
fsm fsm_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
fsm fsm_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
xor_module xor_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
fsm fsm_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
xor_module xor_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
fsm fsm_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
xor_module xor_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
xor_module xor_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
xor_module xor_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
xor_module xor_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
fsm fsm_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
fsm fsm_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
fsm fsm_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
fsm fsm_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
fsm fsm_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
fsm fsm_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
fsm fsm_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
fsm fsm_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
xor_module xor_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
fsm fsm_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
fsm fsm_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
xor_module xor_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
xor_module xor_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
xor_module xor_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
fsm fsm_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
xor_module xor_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
fsm fsm_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
xor_module xor_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
fsm fsm_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
xor_module xor_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
xor_module xor_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
xor_module xor_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
fsm fsm_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
xor_module xor_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
xor_module xor_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
xor_module xor_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
fsm fsm_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
fsm fsm_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
fsm fsm_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
xor_module xor_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
fsm fsm_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
fsm fsm_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
xor_module xor_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
xor_module xor_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
fsm fsm_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
xor_module xor_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
xor_module xor_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
xor_module xor_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
xor_module xor_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
xor_module xor_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
fsm fsm_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
xor_module xor_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
fsm fsm_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
fsm fsm_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
xor_module xor_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
xor_module xor_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
fsm fsm_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
xor_module xor_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
fsm fsm_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
xor_module xor_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
xor_module xor_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
xor_module xor_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
xor_module xor_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
xor_module xor_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
xor_module xor_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
xor_module xor_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
xor_module xor_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
fsm fsm_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
fsm fsm_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
xor_module xor_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
xor_module xor_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
fsm fsm_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
fsm fsm_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
xor_module xor_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
fsm fsm_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
fsm fsm_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
fsm fsm_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
fsm fsm_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
fsm fsm_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
fsm fsm_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
fsm fsm_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
fsm fsm_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
xor_module xor_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
fsm fsm_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
xor_module xor_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
xor_module xor_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
fsm fsm_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
fsm fsm_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
xor_module xor_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
fsm fsm_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
xor_module xor_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
fsm fsm_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
fsm fsm_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
xor_module xor_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
fsm fsm_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
xor_module xor_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
xor_module xor_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
xor_module xor_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
fsm fsm_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
xor_module xor_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
xor_module xor_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
fsm fsm_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
xor_module xor_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
fsm fsm_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
fsm fsm_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
fsm fsm_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
fsm fsm_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
fsm fsm_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
fsm fsm_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
xor_module xor_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
xor_module xor_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
xor_module xor_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
xor_module xor_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
fsm fsm_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
xor_module xor_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
xor_module xor_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
xor_module xor_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
xor_module xor_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
fsm fsm_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
fsm fsm_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
fsm fsm_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
xor_module xor_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
fsm fsm_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
xor_module xor_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
fsm fsm_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
xor_module xor_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
fsm fsm_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
fsm fsm_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
fsm fsm_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
fsm fsm_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
xor_module xor_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
xor_module xor_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
xor_module xor_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
fsm fsm_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
xor_module xor_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
fsm fsm_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
fsm fsm_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
fsm fsm_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
fsm fsm_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
xor_module xor_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
xor_module xor_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
fsm fsm_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
fsm fsm_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
xor_module xor_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
xor_module xor_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
xor_module xor_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
fsm fsm_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
fsm fsm_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
xor_module xor_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
fsm fsm_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
fsm fsm_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
xor_module xor_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
xor_module xor_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
xor_module xor_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
fsm fsm_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
xor_module xor_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
fsm fsm_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
xor_module xor_module_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
fsm fsm_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
fsm fsm_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
fsm fsm_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
fsm fsm_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
fsm fsm_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
fsm fsm_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
xor_module xor_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
xor_module xor_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
xor_module xor_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
fsm fsm_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
fsm fsm_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
xor_module xor_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
xor_module xor_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
xor_module xor_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
xor_module xor_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
fsm fsm_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
xor_module xor_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
fsm fsm_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
xor_module xor_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
fsm fsm_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
xor_module xor_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
fsm fsm_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
xor_module xor_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
xor_module xor_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
fsm fsm_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
xor_module xor_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
xor_module xor_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
fsm fsm_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
fsm fsm_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
xor_module xor_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
fsm fsm_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
xor_module xor_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
xor_module xor_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
xor_module xor_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
xor_module xor_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
fsm fsm_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
xor_module xor_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
fsm fsm_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
fsm fsm_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
fsm fsm_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
xor_module xor_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
xor_module xor_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
fsm fsm_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
xor_module xor_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
fsm fsm_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
xor_module xor_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
fsm fsm_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
xor_module xor_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
fsm fsm_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
fsm fsm_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
fsm fsm_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
fsm fsm_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
xor_module xor_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
fsm fsm_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
xor_module xor_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
xor_module xor_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
fsm fsm_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
fsm fsm_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
xor_module xor_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
fsm fsm_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
fsm fsm_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
fsm fsm_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
fsm fsm_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
fsm fsm_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
xor_module xor_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
xor_module xor_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
fsm fsm_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
fsm fsm_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
xor_module xor_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
fsm fsm_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
xor_module xor_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
xor_module xor_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
fsm fsm_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
fsm fsm_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
xor_module xor_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
xor_module xor_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
xor_module xor_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
xor_module xor_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
fsm fsm_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
xor_module xor_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
xor_module xor_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
xor_module xor_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
fsm fsm_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
xor_module xor_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
xor_module xor_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
xor_module xor_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
xor_module xor_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
fsm fsm_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
fsm fsm_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
fsm fsm_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
xor_module xor_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
xor_module xor_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
fsm fsm_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
fsm fsm_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
xor_module xor_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
xor_module xor_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
xor_module xor_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
xor_module xor_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
fsm fsm_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
xor_module xor_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
xor_module xor_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
fsm fsm_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
xor_module xor_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
fsm fsm_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
fsm fsm_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
fsm fsm_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
fsm fsm_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
xor_module xor_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
fsm fsm_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
fsm fsm_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
fsm fsm_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
fsm fsm_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
fsm fsm_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
xor_module xor_module_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
fsm fsm_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
fsm fsm_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
xor_module xor_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
fsm fsm_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
xor_module xor_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
xor_module xor_module_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
fsm fsm_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
fsm fsm_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
xor_module xor_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
fsm fsm_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
fsm fsm_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
xor_module xor_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
xor_module xor_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
fsm fsm_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
xor_module xor_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
fsm fsm_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
xor_module xor_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
xor_module xor_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
fsm fsm_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
xor_module xor_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
fsm fsm_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
fsm fsm_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
xor_module xor_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
xor_module xor_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
fsm fsm_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
xor_module xor_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
fsm fsm_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
fsm fsm_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
fsm fsm_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
fsm fsm_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
xor_module xor_module_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
xor_module xor_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
fsm fsm_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
xor_module xor_module_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
xor_module xor_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
fsm fsm_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
xor_module xor_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
fsm fsm_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
xor_module xor_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
xor_module xor_module_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
fsm fsm_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
fsm fsm_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
fsm fsm_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
xor_module xor_module_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
fsm fsm_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
xor_module xor_module_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
fsm fsm_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
xor_module xor_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
xor_module xor_module_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
xor_module xor_module_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
fsm fsm_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
xor_module xor_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
fsm fsm_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
fsm fsm_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
xor_module xor_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
xor_module xor_module_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
fsm fsm_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
xor_module xor_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
xor_module xor_module_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
xor_module xor_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
fsm fsm_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
xor_module xor_module_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
fsm fsm_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
xor_module xor_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
fsm fsm_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
xor_module xor_module_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
xor_module xor_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
xor_module xor_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
xor_module xor_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
xor_module xor_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
fsm fsm_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
xor_module xor_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
fsm fsm_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
xor_module xor_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
fsm fsm_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
xor_module xor_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
xor_module xor_module_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
fsm fsm_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
xor_module xor_module_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
fsm fsm_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
fsm fsm_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
fsm fsm_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
xor_module xor_module_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
xor_module xor_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
xor_module xor_module_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
xor_module xor_module_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
fsm fsm_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
fsm fsm_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
xor_module xor_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
fsm fsm_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
fsm fsm_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
xor_module xor_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
xor_module xor_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
xor_module xor_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
xor_module xor_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
fsm fsm_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
xor_module xor_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
fsm fsm_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
fsm fsm_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
fsm fsm_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
xor_module xor_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
xor_module xor_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
fsm fsm_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
xor_module xor_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
xor_module xor_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
fsm fsm_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
fsm fsm_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
fsm fsm_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
reg [619:0]intermediate_reg_2; 
 
fsm fsm_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1239]),.i2(intermediate_reg_1[1238]),.o(intermediate_reg_2[619])); 
xor_module xor_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1237]),.i2(intermediate_reg_1[1236]),.o(intermediate_reg_2[618])); 
fsm fsm_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1235]),.i2(intermediate_reg_1[1234]),.o(intermediate_reg_2[617])); 
xor_module xor_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1233]),.i2(intermediate_reg_1[1232]),.o(intermediate_reg_2[616])); 
xor_module xor_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1231]),.i2(intermediate_reg_1[1230]),.o(intermediate_reg_2[615])); 
fsm fsm_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1229]),.i2(intermediate_reg_1[1228]),.o(intermediate_reg_2[614])); 
fsm fsm_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1227]),.i2(intermediate_reg_1[1226]),.o(intermediate_reg_2[613])); 
fsm fsm_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1225]),.i2(intermediate_reg_1[1224]),.o(intermediate_reg_2[612])); 
fsm fsm_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1223]),.i2(intermediate_reg_1[1222]),.o(intermediate_reg_2[611])); 
xor_module xor_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1221]),.i2(intermediate_reg_1[1220]),.o(intermediate_reg_2[610])); 
fsm fsm_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1219]),.i2(intermediate_reg_1[1218]),.o(intermediate_reg_2[609])); 
xor_module xor_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1217]),.i2(intermediate_reg_1[1216]),.o(intermediate_reg_2[608])); 
fsm fsm_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1215]),.i2(intermediate_reg_1[1214]),.o(intermediate_reg_2[607])); 
fsm fsm_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1213]),.i2(intermediate_reg_1[1212]),.o(intermediate_reg_2[606])); 
xor_module xor_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1211]),.i2(intermediate_reg_1[1210]),.o(intermediate_reg_2[605])); 
xor_module xor_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1209]),.i2(intermediate_reg_1[1208]),.o(intermediate_reg_2[604])); 
fsm fsm_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1207]),.i2(intermediate_reg_1[1206]),.o(intermediate_reg_2[603])); 
fsm fsm_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1205]),.i2(intermediate_reg_1[1204]),.o(intermediate_reg_2[602])); 
xor_module xor_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1203]),.i2(intermediate_reg_1[1202]),.o(intermediate_reg_2[601])); 
xor_module xor_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1201]),.i2(intermediate_reg_1[1200]),.o(intermediate_reg_2[600])); 
fsm fsm_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1199]),.i2(intermediate_reg_1[1198]),.o(intermediate_reg_2[599])); 
fsm fsm_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1197]),.i2(intermediate_reg_1[1196]),.o(intermediate_reg_2[598])); 
xor_module xor_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1195]),.i2(intermediate_reg_1[1194]),.o(intermediate_reg_2[597])); 
fsm fsm_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1193]),.i2(intermediate_reg_1[1192]),.o(intermediate_reg_2[596])); 
fsm fsm_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1191]),.i2(intermediate_reg_1[1190]),.o(intermediate_reg_2[595])); 
fsm fsm_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1189]),.i2(intermediate_reg_1[1188]),.o(intermediate_reg_2[594])); 
xor_module xor_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1187]),.i2(intermediate_reg_1[1186]),.o(intermediate_reg_2[593])); 
fsm fsm_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1185]),.i2(intermediate_reg_1[1184]),.o(intermediate_reg_2[592])); 
fsm fsm_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1183]),.i2(intermediate_reg_1[1182]),.o(intermediate_reg_2[591])); 
fsm fsm_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1181]),.i2(intermediate_reg_1[1180]),.o(intermediate_reg_2[590])); 
fsm fsm_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1179]),.i2(intermediate_reg_1[1178]),.o(intermediate_reg_2[589])); 
fsm fsm_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1177]),.i2(intermediate_reg_1[1176]),.o(intermediate_reg_2[588])); 
xor_module xor_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1175]),.i2(intermediate_reg_1[1174]),.o(intermediate_reg_2[587])); 
xor_module xor_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1173]),.i2(intermediate_reg_1[1172]),.o(intermediate_reg_2[586])); 
fsm fsm_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1171]),.i2(intermediate_reg_1[1170]),.o(intermediate_reg_2[585])); 
fsm fsm_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1169]),.i2(intermediate_reg_1[1168]),.o(intermediate_reg_2[584])); 
fsm fsm_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1167]),.i2(intermediate_reg_1[1166]),.o(intermediate_reg_2[583])); 
fsm fsm_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1165]),.i2(intermediate_reg_1[1164]),.o(intermediate_reg_2[582])); 
fsm fsm_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1163]),.i2(intermediate_reg_1[1162]),.o(intermediate_reg_2[581])); 
xor_module xor_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1161]),.i2(intermediate_reg_1[1160]),.o(intermediate_reg_2[580])); 
xor_module xor_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1159]),.i2(intermediate_reg_1[1158]),.o(intermediate_reg_2[579])); 
xor_module xor_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1157]),.i2(intermediate_reg_1[1156]),.o(intermediate_reg_2[578])); 
xor_module xor_module_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1155]),.i2(intermediate_reg_1[1154]),.o(intermediate_reg_2[577])); 
xor_module xor_module_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1153]),.i2(intermediate_reg_1[1152]),.o(intermediate_reg_2[576])); 
fsm fsm_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1151]),.i2(intermediate_reg_1[1150]),.o(intermediate_reg_2[575])); 
fsm fsm_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1149]),.i2(intermediate_reg_1[1148]),.o(intermediate_reg_2[574])); 
xor_module xor_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1147]),.i2(intermediate_reg_1[1146]),.o(intermediate_reg_2[573])); 
fsm fsm_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1145]),.i2(intermediate_reg_1[1144]),.o(intermediate_reg_2[572])); 
fsm fsm_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1143]),.i2(intermediate_reg_1[1142]),.o(intermediate_reg_2[571])); 
xor_module xor_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1141]),.i2(intermediate_reg_1[1140]),.o(intermediate_reg_2[570])); 
fsm fsm_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1139]),.i2(intermediate_reg_1[1138]),.o(intermediate_reg_2[569])); 
xor_module xor_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1137]),.i2(intermediate_reg_1[1136]),.o(intermediate_reg_2[568])); 
fsm fsm_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1135]),.i2(intermediate_reg_1[1134]),.o(intermediate_reg_2[567])); 
xor_module xor_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1133]),.i2(intermediate_reg_1[1132]),.o(intermediate_reg_2[566])); 
fsm fsm_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1131]),.i2(intermediate_reg_1[1130]),.o(intermediate_reg_2[565])); 
xor_module xor_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1129]),.i2(intermediate_reg_1[1128]),.o(intermediate_reg_2[564])); 
xor_module xor_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1127]),.i2(intermediate_reg_1[1126]),.o(intermediate_reg_2[563])); 
xor_module xor_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1125]),.i2(intermediate_reg_1[1124]),.o(intermediate_reg_2[562])); 
xor_module xor_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1123]),.i2(intermediate_reg_1[1122]),.o(intermediate_reg_2[561])); 
fsm fsm_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1121]),.i2(intermediate_reg_1[1120]),.o(intermediate_reg_2[560])); 
fsm fsm_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1119]),.i2(intermediate_reg_1[1118]),.o(intermediate_reg_2[559])); 
xor_module xor_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1117]),.i2(intermediate_reg_1[1116]),.o(intermediate_reg_2[558])); 
xor_module xor_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1115]),.i2(intermediate_reg_1[1114]),.o(intermediate_reg_2[557])); 
xor_module xor_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1113]),.i2(intermediate_reg_1[1112]),.o(intermediate_reg_2[556])); 
fsm fsm_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1111]),.i2(intermediate_reg_1[1110]),.o(intermediate_reg_2[555])); 
xor_module xor_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1109]),.i2(intermediate_reg_1[1108]),.o(intermediate_reg_2[554])); 
fsm fsm_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1107]),.i2(intermediate_reg_1[1106]),.o(intermediate_reg_2[553])); 
fsm fsm_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1105]),.i2(intermediate_reg_1[1104]),.o(intermediate_reg_2[552])); 
xor_module xor_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1103]),.i2(intermediate_reg_1[1102]),.o(intermediate_reg_2[551])); 
xor_module xor_module_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1101]),.i2(intermediate_reg_1[1100]),.o(intermediate_reg_2[550])); 
xor_module xor_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1099]),.i2(intermediate_reg_1[1098]),.o(intermediate_reg_2[549])); 
fsm fsm_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1097]),.i2(intermediate_reg_1[1096]),.o(intermediate_reg_2[548])); 
xor_module xor_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1095]),.i2(intermediate_reg_1[1094]),.o(intermediate_reg_2[547])); 
xor_module xor_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1093]),.i2(intermediate_reg_1[1092]),.o(intermediate_reg_2[546])); 
fsm fsm_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1091]),.i2(intermediate_reg_1[1090]),.o(intermediate_reg_2[545])); 
fsm fsm_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1089]),.i2(intermediate_reg_1[1088]),.o(intermediate_reg_2[544])); 
xor_module xor_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1087]),.i2(intermediate_reg_1[1086]),.o(intermediate_reg_2[543])); 
xor_module xor_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1085]),.i2(intermediate_reg_1[1084]),.o(intermediate_reg_2[542])); 
xor_module xor_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1083]),.i2(intermediate_reg_1[1082]),.o(intermediate_reg_2[541])); 
fsm fsm_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1081]),.i2(intermediate_reg_1[1080]),.o(intermediate_reg_2[540])); 
xor_module xor_module_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1079]),.i2(intermediate_reg_1[1078]),.o(intermediate_reg_2[539])); 
fsm fsm_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1077]),.i2(intermediate_reg_1[1076]),.o(intermediate_reg_2[538])); 
xor_module xor_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1075]),.i2(intermediate_reg_1[1074]),.o(intermediate_reg_2[537])); 
fsm fsm_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1073]),.i2(intermediate_reg_1[1072]),.o(intermediate_reg_2[536])); 
fsm fsm_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1071]),.i2(intermediate_reg_1[1070]),.o(intermediate_reg_2[535])); 
fsm fsm_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1069]),.i2(intermediate_reg_1[1068]),.o(intermediate_reg_2[534])); 
fsm fsm_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1067]),.i2(intermediate_reg_1[1066]),.o(intermediate_reg_2[533])); 
xor_module xor_module_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1065]),.i2(intermediate_reg_1[1064]),.o(intermediate_reg_2[532])); 
fsm fsm_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1063]),.i2(intermediate_reg_1[1062]),.o(intermediate_reg_2[531])); 
fsm fsm_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1061]),.i2(intermediate_reg_1[1060]),.o(intermediate_reg_2[530])); 
fsm fsm_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1059]),.i2(intermediate_reg_1[1058]),.o(intermediate_reg_2[529])); 
fsm fsm_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1057]),.i2(intermediate_reg_1[1056]),.o(intermediate_reg_2[528])); 
xor_module xor_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1055]),.i2(intermediate_reg_1[1054]),.o(intermediate_reg_2[527])); 
fsm fsm_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1053]),.i2(intermediate_reg_1[1052]),.o(intermediate_reg_2[526])); 
fsm fsm_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1051]),.i2(intermediate_reg_1[1050]),.o(intermediate_reg_2[525])); 
fsm fsm_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1049]),.i2(intermediate_reg_1[1048]),.o(intermediate_reg_2[524])); 
fsm fsm_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1047]),.i2(intermediate_reg_1[1046]),.o(intermediate_reg_2[523])); 
xor_module xor_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1045]),.i2(intermediate_reg_1[1044]),.o(intermediate_reg_2[522])); 
xor_module xor_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1043]),.i2(intermediate_reg_1[1042]),.o(intermediate_reg_2[521])); 
fsm fsm_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1041]),.i2(intermediate_reg_1[1040]),.o(intermediate_reg_2[520])); 
xor_module xor_module_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1039]),.i2(intermediate_reg_1[1038]),.o(intermediate_reg_2[519])); 
fsm fsm_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1037]),.i2(intermediate_reg_1[1036]),.o(intermediate_reg_2[518])); 
fsm fsm_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1035]),.i2(intermediate_reg_1[1034]),.o(intermediate_reg_2[517])); 
xor_module xor_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1033]),.i2(intermediate_reg_1[1032]),.o(intermediate_reg_2[516])); 
fsm fsm_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1031]),.i2(intermediate_reg_1[1030]),.o(intermediate_reg_2[515])); 
fsm fsm_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1029]),.i2(intermediate_reg_1[1028]),.o(intermediate_reg_2[514])); 
xor_module xor_module_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513])); 
fsm fsm_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512])); 
xor_module xor_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511])); 
fsm fsm_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510])); 
xor_module xor_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509])); 
fsm fsm_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508])); 
fsm fsm_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507])); 
xor_module xor_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506])); 
xor_module xor_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505])); 
xor_module xor_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504])); 
fsm fsm_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503])); 
xor_module xor_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502])); 
xor_module xor_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501])); 
fsm fsm_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500])); 
xor_module xor_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499])); 
xor_module xor_module_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498])); 
xor_module xor_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497])); 
fsm fsm_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496])); 
fsm fsm_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495])); 
xor_module xor_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494])); 
fsm fsm_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493])); 
fsm fsm_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492])); 
fsm fsm_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491])); 
fsm fsm_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490])); 
xor_module xor_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489])); 
fsm fsm_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488])); 
fsm fsm_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487])); 
xor_module xor_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486])); 
xor_module xor_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485])); 
fsm fsm_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484])); 
fsm fsm_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483])); 
xor_module xor_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482])); 
xor_module xor_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481])); 
fsm fsm_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480])); 
xor_module xor_module_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
fsm fsm_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478])); 
fsm fsm_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477])); 
xor_module xor_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476])); 
xor_module xor_module_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475])); 
xor_module xor_module_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474])); 
xor_module xor_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473])); 
fsm fsm_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472])); 
fsm fsm_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471])); 
xor_module xor_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470])); 
xor_module xor_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469])); 
fsm fsm_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468])); 
fsm fsm_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467])); 
fsm fsm_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466])); 
xor_module xor_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465])); 
fsm fsm_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464])); 
fsm fsm_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463])); 
fsm fsm_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462])); 
fsm fsm_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461])); 
fsm fsm_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460])); 
xor_module xor_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459])); 
xor_module xor_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458])); 
fsm fsm_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457])); 
fsm fsm_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456])); 
fsm fsm_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455])); 
fsm fsm_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454])); 
xor_module xor_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453])); 
fsm fsm_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452])); 
fsm fsm_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451])); 
xor_module xor_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450])); 
xor_module xor_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449])); 
fsm fsm_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448])); 
xor_module xor_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447])); 
xor_module xor_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446])); 
xor_module xor_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445])); 
xor_module xor_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444])); 
fsm fsm_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443])); 
fsm fsm_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442])); 
xor_module xor_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441])); 
fsm fsm_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440])); 
fsm fsm_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439])); 
fsm fsm_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438])); 
xor_module xor_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437])); 
xor_module xor_module_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436])); 
xor_module xor_module_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435])); 
fsm fsm_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434])); 
fsm fsm_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433])); 
fsm fsm_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432])); 
fsm fsm_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431])); 
xor_module xor_module_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430])); 
xor_module xor_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429])); 
fsm fsm_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428])); 
xor_module xor_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427])); 
fsm fsm_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426])); 
xor_module xor_module_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425])); 
xor_module xor_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424])); 
xor_module xor_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423])); 
xor_module xor_module_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422])); 
fsm fsm_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421])); 
fsm fsm_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420])); 
xor_module xor_module_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419])); 
xor_module xor_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418])); 
fsm fsm_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417])); 
fsm fsm_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416])); 
fsm fsm_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415])); 
xor_module xor_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414])); 
xor_module xor_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413])); 
fsm fsm_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412])); 
fsm fsm_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411])); 
xor_module xor_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410])); 
xor_module xor_module_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409])); 
xor_module xor_module_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408])); 
fsm fsm_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407])); 
fsm fsm_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406])); 
xor_module xor_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405])); 
fsm fsm_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404])); 
xor_module xor_module_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403])); 
fsm fsm_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402])); 
fsm fsm_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401])); 
fsm fsm_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400])); 
xor_module xor_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399])); 
xor_module xor_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398])); 
fsm fsm_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397])); 
xor_module xor_module_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396])); 
fsm fsm_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395])); 
xor_module xor_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394])); 
xor_module xor_module_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393])); 
fsm fsm_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392])); 
xor_module xor_module_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391])); 
xor_module xor_module_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390])); 
xor_module xor_module_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389])); 
xor_module xor_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388])); 
xor_module xor_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387])); 
fsm fsm_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386])); 
fsm fsm_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385])); 
fsm fsm_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384])); 
fsm fsm_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383])); 
fsm fsm_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382])); 
xor_module xor_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
xor_module xor_module_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
xor_module xor_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379])); 
fsm fsm_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378])); 
xor_module xor_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377])); 
xor_module xor_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376])); 
fsm fsm_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375])); 
fsm fsm_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374])); 
xor_module xor_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373])); 
xor_module xor_module_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372])); 
xor_module xor_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371])); 
fsm fsm_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
xor_module xor_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369])); 
xor_module xor_module_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368])); 
fsm fsm_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367])); 
xor_module xor_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366])); 
xor_module xor_module_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365])); 
fsm fsm_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
fsm fsm_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363])); 
xor_module xor_module_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362])); 
xor_module xor_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361])); 
fsm fsm_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360])); 
xor_module xor_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
xor_module xor_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
xor_module xor_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357])); 
fsm fsm_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356])); 
xor_module xor_module_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355])); 
fsm fsm_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354])); 
xor_module xor_module_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353])); 
fsm fsm_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352])); 
xor_module xor_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351])); 
fsm fsm_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350])); 
xor_module xor_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349])); 
fsm fsm_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348])); 
xor_module xor_module_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
fsm fsm_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346])); 
xor_module xor_module_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345])); 
fsm fsm_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
xor_module xor_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343])); 
xor_module xor_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342])); 
xor_module xor_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341])); 
xor_module xor_module_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340])); 
xor_module xor_module_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339])); 
fsm fsm_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338])); 
fsm fsm_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337])); 
xor_module xor_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336])); 
xor_module xor_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
xor_module xor_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334])); 
xor_module xor_module_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333])); 
fsm fsm_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332])); 
fsm fsm_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331])); 
xor_module xor_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
xor_module xor_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
xor_module xor_module_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328])); 
fsm fsm_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
fsm fsm_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326])); 
xor_module xor_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325])); 
xor_module xor_module_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324])); 
fsm fsm_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323])); 
fsm fsm_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322])); 
fsm fsm_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321])); 
xor_module xor_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
xor_module xor_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319])); 
xor_module xor_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318])); 
xor_module xor_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317])); 
fsm fsm_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316])); 
xor_module xor_module_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315])); 
fsm fsm_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314])); 
fsm fsm_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313])); 
xor_module xor_module_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312])); 
xor_module xor_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311])); 
fsm fsm_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310])); 
xor_module xor_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309])); 
xor_module xor_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308])); 
xor_module xor_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307])); 
xor_module xor_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306])); 
fsm fsm_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305])); 
fsm fsm_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304])); 
fsm fsm_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
xor_module xor_module_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302])); 
fsm fsm_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
xor_module xor_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300])); 
xor_module xor_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299])); 
fsm fsm_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298])); 
fsm fsm_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297])); 
xor_module xor_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
xor_module xor_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
fsm fsm_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294])); 
fsm fsm_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
xor_module xor_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292])); 
fsm fsm_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291])); 
xor_module xor_module_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290])); 
xor_module xor_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289])); 
fsm fsm_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288])); 
fsm fsm_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287])); 
xor_module xor_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286])); 
xor_module xor_module_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
xor_module xor_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284])); 
fsm fsm_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
xor_module xor_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282])); 
fsm fsm_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281])); 
xor_module xor_module_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280])); 
xor_module xor_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279])); 
xor_module xor_module_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278])); 
xor_module xor_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277])); 
xor_module xor_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276])); 
fsm fsm_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275])); 
fsm fsm_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
xor_module xor_module_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
xor_module xor_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
fsm fsm_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
xor_module xor_module_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270])); 
fsm fsm_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
xor_module xor_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268])); 
fsm fsm_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267])); 
xor_module xor_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266])); 
fsm fsm_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
xor_module xor_module_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264])); 
fsm fsm_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263])); 
xor_module xor_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
fsm fsm_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261])); 
fsm fsm_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
xor_module xor_module_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259])); 
xor_module xor_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258])); 
fsm fsm_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257])); 
xor_module xor_module_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
fsm fsm_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255])); 
fsm fsm_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254])); 
xor_module xor_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253])); 
xor_module xor_module_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252])); 
xor_module xor_module_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
fsm fsm_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250])); 
fsm fsm_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
xor_module xor_module_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248])); 
xor_module xor_module_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247])); 
fsm fsm_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246])); 
fsm fsm_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
xor_module xor_module_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244])); 
fsm fsm_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243])); 
xor_module xor_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242])); 
xor_module xor_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
fsm fsm_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240])); 
xor_module xor_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239])); 
xor_module xor_module_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
xor_module xor_module_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
fsm fsm_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236])); 
xor_module xor_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235])); 
xor_module xor_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
xor_module xor_module_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233])); 
fsm fsm_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232])); 
xor_module xor_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231])); 
fsm fsm_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230])); 
fsm fsm_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229])); 
fsm fsm_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
fsm fsm_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227])); 
fsm fsm_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
fsm fsm_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
xor_module xor_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224])); 
xor_module xor_module_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223])); 
fsm fsm_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
xor_module xor_module_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221])); 
fsm fsm_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220])); 
xor_module xor_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219])); 
xor_module xor_module_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
xor_module xor_module_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217])); 
xor_module xor_module_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216])); 
xor_module xor_module_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215])); 
fsm fsm_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214])); 
xor_module xor_module_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
xor_module xor_module_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
xor_module xor_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
fsm fsm_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
xor_module xor_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209])); 
fsm fsm_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208])); 
xor_module xor_module_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
fsm fsm_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
xor_module xor_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
xor_module xor_module_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204])); 
xor_module xor_module_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203])); 
xor_module xor_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202])); 
fsm fsm_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201])); 
fsm fsm_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200])); 
fsm fsm_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
xor_module xor_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198])); 
fsm fsm_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197])); 
xor_module xor_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
xor_module xor_module_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195])); 
fsm fsm_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194])); 
fsm fsm_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193])); 
fsm fsm_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
fsm fsm_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
fsm fsm_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190])); 
fsm fsm_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189])); 
fsm fsm_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
fsm fsm_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
fsm fsm_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186])); 
xor_module xor_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185])); 
fsm fsm_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
fsm fsm_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183])); 
fsm fsm_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182])); 
fsm fsm_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181])); 
xor_module xor_module_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180])); 
xor_module xor_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179])); 
xor_module xor_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178])); 
xor_module xor_module_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
xor_module xor_module_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176])); 
fsm fsm_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175])); 
xor_module xor_module_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174])); 
xor_module xor_module_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
fsm fsm_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
xor_module xor_module_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
xor_module xor_module_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
fsm fsm_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169])); 
xor_module xor_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168])); 
fsm fsm_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167])); 
xor_module xor_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166])); 
fsm fsm_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
fsm fsm_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164])); 
fsm fsm_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
xor_module xor_module_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162])); 
xor_module xor_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161])); 
xor_module xor_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160])); 
xor_module xor_module_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
xor_module xor_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158])); 
fsm fsm_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157])); 
xor_module xor_module_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156])); 
xor_module xor_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155])); 
xor_module xor_module_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154])); 
fsm fsm_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153])); 
fsm fsm_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152])); 
xor_module xor_module_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151])); 
xor_module xor_module_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
fsm fsm_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
fsm fsm_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148])); 
xor_module xor_module_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147])); 
fsm fsm_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146])); 
xor_module xor_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145])); 
xor_module xor_module_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144])); 
xor_module xor_module_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143])); 
xor_module xor_module_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142])); 
xor_module xor_module_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141])); 
xor_module xor_module_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140])); 
xor_module xor_module_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139])); 
xor_module xor_module_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138])); 
xor_module xor_module_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
xor_module xor_module_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136])); 
fsm fsm_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135])); 
fsm fsm_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
xor_module xor_module_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133])); 
fsm fsm_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132])); 
xor_module xor_module_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131])); 
fsm fsm_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130])); 
xor_module xor_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129])); 
fsm fsm_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
xor_module xor_module_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
fsm fsm_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126])); 
fsm fsm_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
fsm fsm_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124])); 
xor_module xor_module_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123])); 
xor_module xor_module_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
xor_module xor_module_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121])); 
fsm fsm_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120])); 
xor_module xor_module_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119])); 
xor_module xor_module_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118])); 
fsm fsm_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117])); 
fsm fsm_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116])); 
fsm fsm_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115])); 
xor_module xor_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
xor_module xor_module_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113])); 
fsm fsm_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
xor_module xor_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111])); 
xor_module xor_module_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
xor_module xor_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
xor_module xor_module_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
xor_module xor_module_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107])); 
xor_module xor_module_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
fsm fsm_inst_2_514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105])); 
xor_module xor_module_inst_2_515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104])); 
xor_module xor_module_inst_2_516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
fsm fsm_inst_2_517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102])); 
fsm fsm_inst_2_518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
xor_module xor_module_inst_2_519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100])); 
fsm fsm_inst_2_520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99])); 
fsm fsm_inst_2_521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98])); 
fsm fsm_inst_2_522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
xor_module xor_module_inst_2_523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96])); 
xor_module xor_module_inst_2_524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95])); 
fsm fsm_inst_2_525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94])); 
fsm fsm_inst_2_526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
xor_module xor_module_inst_2_527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92])); 
xor_module xor_module_inst_2_528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91])); 
xor_module xor_module_inst_2_529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
fsm fsm_inst_2_530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89])); 
fsm fsm_inst_2_531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88])); 
fsm fsm_inst_2_532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
fsm fsm_inst_2_533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
xor_module xor_module_inst_2_534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
xor_module xor_module_inst_2_535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
fsm fsm_inst_2_536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
fsm fsm_inst_2_537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82])); 
fsm fsm_inst_2_538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
fsm fsm_inst_2_539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80])); 
fsm fsm_inst_2_540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79])); 
fsm fsm_inst_2_541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78])); 
fsm fsm_inst_2_542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
fsm fsm_inst_2_543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76])); 
fsm fsm_inst_2_544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
xor_module xor_module_inst_2_545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74])); 
fsm fsm_inst_2_546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73])); 
fsm fsm_inst_2_547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72])); 
fsm fsm_inst_2_548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71])); 
xor_module xor_module_inst_2_549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
fsm fsm_inst_2_550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69])); 
fsm fsm_inst_2_551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68])); 
fsm fsm_inst_2_552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67])); 
fsm fsm_inst_2_553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66])); 
xor_module xor_module_inst_2_554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65])); 
fsm fsm_inst_2_555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64])); 
fsm fsm_inst_2_556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
fsm fsm_inst_2_557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
xor_module xor_module_inst_2_558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
fsm fsm_inst_2_559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60])); 
xor_module xor_module_inst_2_560(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59])); 
fsm fsm_inst_2_561(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
fsm fsm_inst_2_562(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57])); 
xor_module xor_module_inst_2_563(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56])); 
xor_module xor_module_inst_2_564(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55])); 
xor_module xor_module_inst_2_565(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54])); 
fsm fsm_inst_2_566(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
fsm fsm_inst_2_567(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
fsm fsm_inst_2_568(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51])); 
fsm fsm_inst_2_569(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
xor_module xor_module_inst_2_570(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
fsm fsm_inst_2_571(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48])); 
fsm fsm_inst_2_572(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47])); 
fsm fsm_inst_2_573(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46])); 
fsm fsm_inst_2_574(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45])); 
fsm fsm_inst_2_575(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44])); 
xor_module xor_module_inst_2_576(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
fsm fsm_inst_2_577(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42])); 
fsm fsm_inst_2_578(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
xor_module xor_module_inst_2_579(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40])); 
xor_module xor_module_inst_2_580(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39])); 
xor_module xor_module_inst_2_581(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38])); 
fsm fsm_inst_2_582(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
fsm fsm_inst_2_583(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36])); 
fsm fsm_inst_2_584(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35])); 
fsm fsm_inst_2_585(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34])); 
xor_module xor_module_inst_2_586(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33])); 
fsm fsm_inst_2_587(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32])); 
fsm fsm_inst_2_588(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
xor_module xor_module_inst_2_589(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
xor_module xor_module_inst_2_590(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29])); 
fsm fsm_inst_2_591(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
fsm fsm_inst_2_592(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27])); 
xor_module xor_module_inst_2_593(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26])); 
xor_module xor_module_inst_2_594(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25])); 
xor_module xor_module_inst_2_595(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
xor_module xor_module_inst_2_596(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23])); 
xor_module xor_module_inst_2_597(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22])); 
xor_module xor_module_inst_2_598(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21])); 
xor_module xor_module_inst_2_599(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20])); 
fsm fsm_inst_2_600(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
fsm fsm_inst_2_601(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18])); 
xor_module xor_module_inst_2_602(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17])); 
xor_module xor_module_inst_2_603(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
xor_module xor_module_inst_2_604(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15])); 
fsm fsm_inst_2_605(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14])); 
xor_module xor_module_inst_2_606(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13])); 
fsm fsm_inst_2_607(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12])); 
xor_module xor_module_inst_2_608(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11])); 
fsm fsm_inst_2_609(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10])); 
fsm fsm_inst_2_610(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
xor_module xor_module_inst_2_611(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8])); 
xor_module xor_module_inst_2_612(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
xor_module xor_module_inst_2_613(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6])); 
xor_module xor_module_inst_2_614(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5])); 
xor_module xor_module_inst_2_615(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
xor_module xor_module_inst_2_616(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
fsm fsm_inst_2_617(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2])); 
xor_module xor_module_inst_2_618(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
fsm fsm_inst_2_619(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0])); 
always@(posedge clk) begin 
outp [619:0] <= intermediate_reg_2; 
outp[1059:620] <= intermediate_reg_2[439:0] ; 
end 
endmodule 
 

module interface_11(input [1595:0] inp, output reg [171:0] outp, input clk, input reset);
reg [1595:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [797:0]intermediate_reg_1; 
 
xor_module xor_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
fsm fsm_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
xor_module xor_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
xor_module xor_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
xor_module xor_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
fsm fsm_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
xor_module xor_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
xor_module xor_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
xor_module xor_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
xor_module xor_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
fsm fsm_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
fsm fsm_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
xor_module xor_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
xor_module xor_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
xor_module xor_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
fsm fsm_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
fsm fsm_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
xor_module xor_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
fsm fsm_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
xor_module xor_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
fsm fsm_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
xor_module xor_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
xor_module xor_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
xor_module xor_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
xor_module xor_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
fsm fsm_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
xor_module xor_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
xor_module xor_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
xor_module xor_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
fsm fsm_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
fsm fsm_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
fsm fsm_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
fsm fsm_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
fsm fsm_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
xor_module xor_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
fsm fsm_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
fsm fsm_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
xor_module xor_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
xor_module xor_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
xor_module xor_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
fsm fsm_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
xor_module xor_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
xor_module xor_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
fsm fsm_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
xor_module xor_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
fsm fsm_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
fsm fsm_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
xor_module xor_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
fsm fsm_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
fsm fsm_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
fsm fsm_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
fsm fsm_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
xor_module xor_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
xor_module xor_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
fsm fsm_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687])); 
xor_module xor_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
fsm fsm_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
xor_module xor_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
fsm fsm_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
xor_module xor_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
fsm fsm_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
xor_module xor_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
fsm fsm_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
fsm fsm_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
xor_module xor_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
fsm fsm_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
fsm fsm_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
fsm fsm_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
fsm fsm_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
xor_module xor_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
fsm fsm_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
fsm fsm_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
fsm fsm_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
xor_module xor_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
xor_module xor_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
xor_module xor_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
fsm fsm_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
xor_module xor_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
fsm fsm_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
fsm fsm_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
fsm fsm_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640])); 
fsm fsm_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
fsm fsm_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
xor_module xor_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
xor_module xor_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
fsm fsm_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
fsm fsm_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
fsm fsm_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
xor_module xor_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
fsm fsm_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
fsm fsm_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
xor_module xor_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
xor_module xor_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
xor_module xor_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
fsm fsm_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
fsm fsm_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
xor_module xor_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
fsm fsm_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
fsm fsm_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
fsm fsm_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
fsm fsm_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
fsm fsm_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
xor_module xor_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
fsm fsm_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
xor_module xor_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
xor_module xor_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
xor_module xor_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
fsm fsm_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
fsm fsm_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
xor_module xor_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
fsm fsm_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
fsm fsm_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
fsm fsm_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
fsm fsm_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
fsm fsm_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
fsm fsm_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
fsm fsm_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
fsm fsm_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
xor_module xor_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
fsm fsm_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
xor_module xor_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
fsm fsm_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
xor_module xor_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
xor_module xor_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
xor_module xor_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
xor_module xor_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
xor_module xor_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
xor_module xor_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
fsm fsm_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
xor_module xor_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
fsm fsm_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
fsm fsm_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
fsm fsm_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
xor_module xor_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
xor_module xor_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
fsm fsm_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
xor_module xor_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
fsm fsm_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
xor_module xor_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
xor_module xor_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
fsm fsm_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
xor_module xor_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
xor_module xor_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
fsm fsm_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
fsm fsm_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
xor_module xor_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
fsm fsm_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
fsm fsm_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
fsm fsm_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
fsm fsm_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
xor_module xor_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
fsm fsm_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
fsm fsm_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
fsm fsm_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
fsm fsm_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
fsm fsm_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
fsm fsm_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
fsm fsm_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
fsm fsm_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
fsm fsm_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
fsm fsm_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
fsm fsm_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
fsm fsm_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
xor_module xor_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
fsm fsm_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
fsm fsm_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
xor_module xor_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
xor_module xor_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
fsm fsm_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
fsm fsm_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
xor_module xor_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
xor_module xor_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
fsm fsm_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
fsm fsm_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
xor_module xor_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
fsm fsm_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
fsm fsm_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
fsm fsm_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
fsm fsm_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
fsm fsm_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
xor_module xor_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
fsm fsm_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
fsm fsm_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
xor_module xor_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
fsm fsm_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
fsm fsm_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
xor_module xor_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
fsm fsm_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
fsm fsm_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
fsm fsm_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
xor_module xor_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
fsm fsm_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
fsm fsm_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
fsm fsm_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
fsm fsm_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
fsm fsm_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
fsm fsm_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
fsm fsm_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
xor_module xor_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
fsm fsm_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
xor_module xor_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
xor_module xor_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
fsm fsm_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
fsm fsm_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
xor_module xor_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
fsm fsm_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
xor_module xor_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
fsm fsm_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
xor_module xor_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
fsm fsm_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
fsm fsm_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
fsm fsm_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
fsm fsm_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
fsm fsm_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
xor_module xor_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
fsm fsm_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
fsm fsm_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
fsm fsm_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
xor_module xor_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
fsm fsm_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
xor_module xor_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
fsm fsm_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
xor_module xor_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
fsm fsm_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
fsm fsm_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
xor_module xor_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
fsm fsm_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
fsm fsm_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
fsm fsm_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
fsm fsm_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
fsm fsm_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
fsm fsm_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
fsm fsm_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
fsm fsm_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
xor_module xor_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
fsm fsm_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
xor_module xor_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
fsm fsm_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
fsm fsm_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
fsm fsm_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
xor_module xor_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
fsm fsm_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
fsm fsm_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
xor_module xor_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
fsm fsm_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
fsm fsm_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
fsm fsm_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
fsm fsm_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
fsm fsm_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
fsm fsm_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
fsm fsm_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
fsm fsm_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
fsm fsm_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
fsm fsm_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
fsm fsm_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
xor_module xor_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
xor_module xor_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
fsm fsm_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
xor_module xor_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
xor_module xor_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
fsm fsm_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
fsm fsm_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
xor_module xor_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
fsm fsm_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
fsm fsm_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
fsm fsm_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
fsm fsm_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
fsm fsm_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
fsm fsm_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
fsm fsm_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
fsm fsm_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
xor_module xor_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
fsm fsm_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
xor_module xor_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
fsm fsm_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
fsm fsm_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
fsm fsm_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
fsm fsm_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
xor_module xor_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
fsm fsm_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
fsm fsm_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
fsm fsm_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
xor_module xor_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
xor_module xor_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
xor_module xor_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
fsm fsm_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
fsm fsm_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
xor_module xor_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
xor_module xor_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
xor_module xor_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
fsm fsm_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
xor_module xor_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
xor_module xor_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
xor_module xor_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
fsm fsm_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
xor_module xor_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
fsm fsm_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
fsm fsm_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
fsm fsm_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
fsm fsm_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
fsm fsm_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
fsm fsm_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
fsm fsm_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
fsm fsm_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
fsm fsm_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
xor_module xor_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
fsm fsm_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
fsm fsm_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
fsm fsm_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
fsm fsm_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
xor_module xor_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
xor_module xor_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
fsm fsm_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
xor_module xor_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
fsm fsm_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
xor_module xor_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
xor_module xor_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
fsm fsm_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
xor_module xor_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
xor_module xor_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
fsm fsm_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
xor_module xor_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
xor_module xor_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
xor_module xor_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
fsm fsm_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
fsm fsm_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
xor_module xor_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
xor_module xor_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
xor_module xor_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
fsm fsm_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
xor_module xor_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
fsm fsm_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
fsm fsm_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
fsm fsm_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
fsm fsm_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
fsm fsm_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
fsm fsm_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
fsm fsm_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
xor_module xor_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
xor_module xor_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
fsm fsm_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
fsm fsm_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
fsm fsm_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
xor_module xor_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
fsm fsm_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
xor_module xor_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
xor_module xor_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
fsm fsm_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
fsm fsm_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
xor_module xor_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
xor_module xor_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
xor_module xor_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
fsm fsm_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
xor_module xor_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
fsm fsm_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
fsm fsm_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
fsm fsm_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
xor_module xor_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
xor_module xor_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
fsm fsm_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
fsm fsm_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
xor_module xor_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
xor_module xor_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
fsm fsm_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
xor_module xor_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
xor_module xor_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
fsm fsm_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
xor_module xor_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
fsm fsm_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
fsm fsm_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
xor_module xor_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
fsm fsm_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
fsm fsm_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
fsm fsm_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
xor_module xor_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
fsm fsm_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
fsm fsm_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
xor_module xor_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
fsm fsm_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
fsm fsm_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
xor_module xor_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
xor_module xor_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
fsm fsm_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
fsm fsm_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
fsm fsm_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
xor_module xor_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
fsm fsm_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
fsm fsm_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
fsm fsm_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
xor_module xor_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
xor_module xor_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
fsm fsm_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
fsm fsm_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
fsm fsm_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
xor_module xor_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
xor_module xor_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
fsm fsm_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
fsm fsm_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
xor_module xor_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
fsm fsm_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
xor_module xor_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
fsm fsm_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
xor_module xor_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
fsm fsm_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
fsm fsm_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
xor_module xor_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
fsm fsm_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
xor_module xor_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
fsm fsm_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
fsm fsm_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
fsm fsm_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
xor_module xor_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
fsm fsm_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
xor_module xor_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
xor_module xor_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
xor_module xor_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
fsm fsm_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
fsm fsm_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
fsm fsm_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
fsm fsm_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
xor_module xor_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
fsm fsm_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
xor_module xor_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
xor_module xor_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
fsm fsm_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
fsm fsm_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
fsm fsm_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
fsm fsm_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
fsm fsm_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
fsm fsm_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
fsm fsm_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
xor_module xor_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
fsm fsm_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
fsm fsm_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
xor_module xor_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
fsm fsm_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
fsm fsm_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
fsm fsm_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
xor_module xor_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
xor_module xor_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
xor_module xor_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
xor_module xor_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
fsm fsm_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
xor_module xor_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
fsm fsm_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
fsm fsm_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
xor_module xor_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
xor_module xor_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
xor_module xor_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
xor_module xor_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
xor_module xor_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
fsm fsm_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
xor_module xor_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
fsm fsm_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
fsm fsm_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
reg [398:0]intermediate_reg_2; 
 
xor_module xor_module_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398])); 
fsm fsm_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397])); 
xor_module xor_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396])); 
fsm fsm_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395])); 
fsm fsm_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394])); 
fsm fsm_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393])); 
xor_module xor_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392])); 
xor_module xor_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391])); 
fsm fsm_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390])); 
xor_module xor_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389])); 
fsm fsm_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388])); 
xor_module xor_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387])); 
xor_module xor_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386])); 
xor_module xor_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385])); 
xor_module xor_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384])); 
fsm fsm_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383])); 
fsm fsm_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382])); 
xor_module xor_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
fsm fsm_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
xor_module xor_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379])); 
fsm fsm_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378])); 
xor_module xor_module_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377])); 
fsm fsm_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376])); 
xor_module xor_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375])); 
xor_module xor_module_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374])); 
fsm fsm_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373])); 
fsm fsm_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372])); 
fsm fsm_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371])); 
fsm fsm_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
fsm fsm_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369])); 
xor_module xor_module_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368])); 
xor_module xor_module_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367])); 
xor_module xor_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366])); 
xor_module xor_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365])); 
fsm fsm_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
xor_module xor_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363])); 
fsm fsm_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362])); 
xor_module xor_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361])); 
xor_module xor_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360])); 
fsm fsm_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
fsm fsm_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
xor_module xor_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357])); 
fsm fsm_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356])); 
fsm fsm_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355])); 
xor_module xor_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354])); 
xor_module xor_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353])); 
xor_module xor_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352])); 
xor_module xor_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351])); 
fsm fsm_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350])); 
xor_module xor_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349])); 
xor_module xor_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348])); 
xor_module xor_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
xor_module xor_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346])); 
fsm fsm_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345])); 
xor_module xor_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
fsm fsm_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343])); 
xor_module xor_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342])); 
fsm fsm_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341])); 
fsm fsm_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340])); 
xor_module xor_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339])); 
fsm fsm_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338])); 
fsm fsm_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337])); 
fsm fsm_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336])); 
fsm fsm_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
fsm fsm_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334])); 
fsm fsm_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333])); 
fsm fsm_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332])); 
xor_module xor_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331])); 
fsm fsm_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
fsm fsm_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
fsm fsm_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328])); 
xor_module xor_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
fsm fsm_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326])); 
xor_module xor_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325])); 
xor_module xor_module_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324])); 
xor_module xor_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323])); 
fsm fsm_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322])); 
xor_module xor_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321])); 
fsm fsm_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
xor_module xor_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319])); 
fsm fsm_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318])); 
fsm fsm_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317])); 
xor_module xor_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316])); 
fsm fsm_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315])); 
xor_module xor_module_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314])); 
fsm fsm_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313])); 
xor_module xor_module_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312])); 
fsm fsm_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311])); 
xor_module xor_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310])); 
fsm fsm_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309])); 
xor_module xor_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308])); 
xor_module xor_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307])); 
xor_module xor_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306])); 
xor_module xor_module_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305])); 
xor_module xor_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304])); 
fsm fsm_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
xor_module xor_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302])); 
fsm fsm_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
xor_module xor_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300])); 
xor_module xor_module_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299])); 
fsm fsm_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298])); 
xor_module xor_module_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297])); 
fsm fsm_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
xor_module xor_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
xor_module xor_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294])); 
xor_module xor_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
fsm fsm_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292])); 
fsm fsm_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291])); 
xor_module xor_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290])); 
xor_module xor_module_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289])); 
fsm fsm_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288])); 
xor_module xor_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287])); 
fsm fsm_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286])); 
fsm fsm_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
xor_module xor_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284])); 
xor_module xor_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
xor_module xor_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282])); 
xor_module xor_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281])); 
xor_module xor_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280])); 
xor_module xor_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279])); 
xor_module xor_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278])); 
fsm fsm_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277])); 
fsm fsm_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276])); 
xor_module xor_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275])); 
fsm fsm_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
fsm fsm_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
xor_module xor_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
xor_module xor_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
fsm fsm_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270])); 
fsm fsm_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
xor_module xor_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268])); 
xor_module xor_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267])); 
xor_module xor_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266])); 
xor_module xor_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
xor_module xor_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264])); 
fsm fsm_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263])); 
xor_module xor_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
fsm fsm_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261])); 
xor_module xor_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
xor_module xor_module_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259])); 
fsm fsm_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258])); 
xor_module xor_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257])); 
xor_module xor_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
xor_module xor_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255])); 
fsm fsm_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254])); 
fsm fsm_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253])); 
xor_module xor_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252])); 
fsm fsm_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
xor_module xor_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250])); 
xor_module xor_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
fsm fsm_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248])); 
fsm fsm_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247])); 
xor_module xor_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246])); 
fsm fsm_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
xor_module xor_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244])); 
xor_module xor_module_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243])); 
fsm fsm_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242])); 
xor_module xor_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
fsm fsm_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240])); 
xor_module xor_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239])); 
xor_module xor_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
xor_module xor_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
xor_module xor_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236])); 
xor_module xor_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235])); 
xor_module xor_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
fsm fsm_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233])); 
xor_module xor_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232])); 
fsm fsm_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231])); 
fsm fsm_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230])); 
fsm fsm_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229])); 
fsm fsm_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
fsm fsm_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227])); 
xor_module xor_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
xor_module xor_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
fsm fsm_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224])); 
xor_module xor_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223])); 
xor_module xor_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
xor_module xor_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221])); 
xor_module xor_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220])); 
xor_module xor_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219])); 
fsm fsm_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
fsm fsm_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217])); 
fsm fsm_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216])); 
fsm fsm_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215])); 
xor_module xor_module_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214])); 
fsm fsm_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
xor_module xor_module_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
fsm fsm_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
fsm fsm_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
fsm fsm_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209])); 
xor_module xor_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208])); 
fsm fsm_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
xor_module xor_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
xor_module xor_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
xor_module xor_module_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204])); 
xor_module xor_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203])); 
fsm fsm_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202])); 
fsm fsm_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201])); 
xor_module xor_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200])); 
fsm fsm_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
fsm fsm_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198])); 
fsm fsm_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197])); 
fsm fsm_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
xor_module xor_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195])); 
fsm fsm_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194])); 
xor_module xor_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193])); 
xor_module xor_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
xor_module xor_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
xor_module xor_module_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190])); 
fsm fsm_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189])); 
xor_module xor_module_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
fsm fsm_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
xor_module xor_module_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186])); 
xor_module xor_module_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185])); 
xor_module xor_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
fsm fsm_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183])); 
fsm fsm_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182])); 
fsm fsm_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181])); 
fsm fsm_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180])); 
fsm fsm_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179])); 
xor_module xor_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178])); 
xor_module xor_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
fsm fsm_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176])); 
xor_module xor_module_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175])); 
fsm fsm_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174])); 
xor_module xor_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
fsm fsm_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
fsm fsm_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
xor_module xor_module_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
xor_module xor_module_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169])); 
xor_module xor_module_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168])); 
fsm fsm_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167])); 
xor_module xor_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166])); 
xor_module xor_module_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
xor_module xor_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164])); 
xor_module xor_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
fsm fsm_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162])); 
fsm fsm_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161])); 
xor_module xor_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160])); 
fsm fsm_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
xor_module xor_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158])); 
fsm fsm_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157])); 
xor_module xor_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156])); 
fsm fsm_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155])); 
xor_module xor_module_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154])); 
xor_module xor_module_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153])); 
fsm fsm_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152])); 
fsm fsm_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151])); 
fsm fsm_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
fsm fsm_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
fsm fsm_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148])); 
fsm fsm_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147])); 
xor_module xor_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146])); 
fsm fsm_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145])); 
fsm fsm_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144])); 
xor_module xor_module_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143])); 
fsm fsm_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142])); 
fsm fsm_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141])); 
fsm fsm_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140])); 
fsm fsm_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139])); 
fsm fsm_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138])); 
xor_module xor_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
xor_module xor_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136])); 
fsm fsm_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135])); 
fsm fsm_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
xor_module xor_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133])); 
xor_module xor_module_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132])); 
fsm fsm_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131])); 
xor_module xor_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130])); 
fsm fsm_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129])); 
fsm fsm_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
fsm fsm_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
fsm fsm_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126])); 
xor_module xor_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
fsm fsm_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124])); 
fsm fsm_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123])); 
xor_module xor_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
xor_module xor_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121])); 
fsm fsm_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120])); 
fsm fsm_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119])); 
xor_module xor_module_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118])); 
fsm fsm_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117])); 
xor_module xor_module_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116])); 
xor_module xor_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115])); 
xor_module xor_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
xor_module xor_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113])); 
xor_module xor_module_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
xor_module xor_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111])); 
fsm fsm_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
xor_module xor_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
fsm fsm_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
xor_module xor_module_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107])); 
fsm fsm_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
xor_module xor_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105])); 
fsm fsm_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104])); 
fsm fsm_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
fsm fsm_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102])); 
fsm fsm_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
fsm fsm_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100])); 
xor_module xor_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99])); 
xor_module xor_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98])); 
xor_module xor_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
fsm fsm_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96])); 
fsm fsm_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95])); 
fsm fsm_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94])); 
xor_module xor_module_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
fsm fsm_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92])); 
xor_module xor_module_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91])); 
xor_module xor_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
fsm fsm_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89])); 
xor_module xor_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88])); 
xor_module xor_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
xor_module xor_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
xor_module xor_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
xor_module xor_module_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
xor_module xor_module_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
xor_module xor_module_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82])); 
fsm fsm_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
fsm fsm_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80])); 
xor_module xor_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79])); 
fsm fsm_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78])); 
fsm fsm_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
xor_module xor_module_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76])); 
xor_module xor_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
xor_module xor_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74])); 
xor_module xor_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73])); 
fsm fsm_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72])); 
xor_module xor_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71])); 
xor_module xor_module_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
fsm fsm_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69])); 
fsm fsm_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68])); 
fsm fsm_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67])); 
fsm fsm_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66])); 
xor_module xor_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65])); 
fsm fsm_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64])); 
xor_module xor_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
xor_module xor_module_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
fsm fsm_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
xor_module xor_module_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60])); 
fsm fsm_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59])); 
xor_module xor_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
fsm fsm_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57])); 
fsm fsm_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56])); 
xor_module xor_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55])); 
fsm fsm_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54])); 
fsm fsm_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
fsm fsm_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
fsm fsm_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51])); 
fsm fsm_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
xor_module xor_module_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
fsm fsm_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48])); 
xor_module xor_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47])); 
fsm fsm_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46])); 
xor_module xor_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45])); 
xor_module xor_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44])); 
fsm fsm_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
fsm fsm_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42])); 
xor_module xor_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
fsm fsm_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40])); 
fsm fsm_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39])); 
fsm fsm_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38])); 
xor_module xor_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
xor_module xor_module_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36])); 
fsm fsm_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35])); 
xor_module xor_module_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34])); 
fsm fsm_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33])); 
xor_module xor_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32])); 
fsm fsm_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
fsm fsm_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
fsm fsm_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29])); 
fsm fsm_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
xor_module xor_module_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27])); 
fsm fsm_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26])); 
fsm fsm_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25])); 
fsm fsm_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
fsm fsm_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23])); 
fsm fsm_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22])); 
fsm fsm_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21])); 
fsm fsm_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20])); 
xor_module xor_module_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
fsm fsm_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18])); 
fsm fsm_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17])); 
fsm fsm_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
xor_module xor_module_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15])); 
xor_module xor_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14])); 
xor_module xor_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13])); 
fsm fsm_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12])); 
fsm fsm_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11])); 
xor_module xor_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10])); 
fsm fsm_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
xor_module xor_module_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8])); 
xor_module xor_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
xor_module xor_module_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6])); 
xor_module xor_module_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5])); 
fsm fsm_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
xor_module xor_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
xor_module xor_module_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2])); 
fsm fsm_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
fsm fsm_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0])); 
wire [397:0]intermediate_wire_3; 
assign intermediate_wire_3[397] = intermediate_reg_2[398]^intermediate_reg_2[397] ; 
assign intermediate_wire_3[396:0] = intermediate_reg_2[396:0] ; 
reg [198:0]intermediate_reg_3; 
 
xor_module xor_module_inst_3_0(.clk(clk),.reset(reset),.i1(intermediate_wire_3[397]),.i2(intermediate_wire_3[396]),.o(intermediate_reg_3[198])); 
fsm fsm_inst_3_1(.clk(clk),.reset(reset),.i1(intermediate_wire_3[395]),.i2(intermediate_wire_3[394]),.o(intermediate_reg_3[197])); 
fsm fsm_inst_3_2(.clk(clk),.reset(reset),.i1(intermediate_wire_3[393]),.i2(intermediate_wire_3[392]),.o(intermediate_reg_3[196])); 
fsm fsm_inst_3_3(.clk(clk),.reset(reset),.i1(intermediate_wire_3[391]),.i2(intermediate_wire_3[390]),.o(intermediate_reg_3[195])); 
xor_module xor_module_inst_3_4(.clk(clk),.reset(reset),.i1(intermediate_wire_3[389]),.i2(intermediate_wire_3[388]),.o(intermediate_reg_3[194])); 
xor_module xor_module_inst_3_5(.clk(clk),.reset(reset),.i1(intermediate_wire_3[387]),.i2(intermediate_wire_3[386]),.o(intermediate_reg_3[193])); 
xor_module xor_module_inst_3_6(.clk(clk),.reset(reset),.i1(intermediate_wire_3[385]),.i2(intermediate_wire_3[384]),.o(intermediate_reg_3[192])); 
xor_module xor_module_inst_3_7(.clk(clk),.reset(reset),.i1(intermediate_wire_3[383]),.i2(intermediate_wire_3[382]),.o(intermediate_reg_3[191])); 
fsm fsm_inst_3_8(.clk(clk),.reset(reset),.i1(intermediate_wire_3[381]),.i2(intermediate_wire_3[380]),.o(intermediate_reg_3[190])); 
fsm fsm_inst_3_9(.clk(clk),.reset(reset),.i1(intermediate_wire_3[379]),.i2(intermediate_wire_3[378]),.o(intermediate_reg_3[189])); 
xor_module xor_module_inst_3_10(.clk(clk),.reset(reset),.i1(intermediate_wire_3[377]),.i2(intermediate_wire_3[376]),.o(intermediate_reg_3[188])); 
fsm fsm_inst_3_11(.clk(clk),.reset(reset),.i1(intermediate_wire_3[375]),.i2(intermediate_wire_3[374]),.o(intermediate_reg_3[187])); 
fsm fsm_inst_3_12(.clk(clk),.reset(reset),.i1(intermediate_wire_3[373]),.i2(intermediate_wire_3[372]),.o(intermediate_reg_3[186])); 
fsm fsm_inst_3_13(.clk(clk),.reset(reset),.i1(intermediate_wire_3[371]),.i2(intermediate_wire_3[370]),.o(intermediate_reg_3[185])); 
fsm fsm_inst_3_14(.clk(clk),.reset(reset),.i1(intermediate_wire_3[369]),.i2(intermediate_wire_3[368]),.o(intermediate_reg_3[184])); 
fsm fsm_inst_3_15(.clk(clk),.reset(reset),.i1(intermediate_wire_3[367]),.i2(intermediate_wire_3[366]),.o(intermediate_reg_3[183])); 
fsm fsm_inst_3_16(.clk(clk),.reset(reset),.i1(intermediate_wire_3[365]),.i2(intermediate_wire_3[364]),.o(intermediate_reg_3[182])); 
fsm fsm_inst_3_17(.clk(clk),.reset(reset),.i1(intermediate_wire_3[363]),.i2(intermediate_wire_3[362]),.o(intermediate_reg_3[181])); 
fsm fsm_inst_3_18(.clk(clk),.reset(reset),.i1(intermediate_wire_3[361]),.i2(intermediate_wire_3[360]),.o(intermediate_reg_3[180])); 
fsm fsm_inst_3_19(.clk(clk),.reset(reset),.i1(intermediate_wire_3[359]),.i2(intermediate_wire_3[358]),.o(intermediate_reg_3[179])); 
fsm fsm_inst_3_20(.clk(clk),.reset(reset),.i1(intermediate_wire_3[357]),.i2(intermediate_wire_3[356]),.o(intermediate_reg_3[178])); 
xor_module xor_module_inst_3_21(.clk(clk),.reset(reset),.i1(intermediate_wire_3[355]),.i2(intermediate_wire_3[354]),.o(intermediate_reg_3[177])); 
xor_module xor_module_inst_3_22(.clk(clk),.reset(reset),.i1(intermediate_wire_3[353]),.i2(intermediate_wire_3[352]),.o(intermediate_reg_3[176])); 
fsm fsm_inst_3_23(.clk(clk),.reset(reset),.i1(intermediate_wire_3[351]),.i2(intermediate_wire_3[350]),.o(intermediate_reg_3[175])); 
fsm fsm_inst_3_24(.clk(clk),.reset(reset),.i1(intermediate_wire_3[349]),.i2(intermediate_wire_3[348]),.o(intermediate_reg_3[174])); 
fsm fsm_inst_3_25(.clk(clk),.reset(reset),.i1(intermediate_wire_3[347]),.i2(intermediate_wire_3[346]),.o(intermediate_reg_3[173])); 
xor_module xor_module_inst_3_26(.clk(clk),.reset(reset),.i1(intermediate_wire_3[345]),.i2(intermediate_wire_3[344]),.o(intermediate_reg_3[172])); 
fsm fsm_inst_3_27(.clk(clk),.reset(reset),.i1(intermediate_wire_3[343]),.i2(intermediate_wire_3[342]),.o(intermediate_reg_3[171])); 
xor_module xor_module_inst_3_28(.clk(clk),.reset(reset),.i1(intermediate_wire_3[341]),.i2(intermediate_wire_3[340]),.o(intermediate_reg_3[170])); 
fsm fsm_inst_3_29(.clk(clk),.reset(reset),.i1(intermediate_wire_3[339]),.i2(intermediate_wire_3[338]),.o(intermediate_reg_3[169])); 
xor_module xor_module_inst_3_30(.clk(clk),.reset(reset),.i1(intermediate_wire_3[337]),.i2(intermediate_wire_3[336]),.o(intermediate_reg_3[168])); 
xor_module xor_module_inst_3_31(.clk(clk),.reset(reset),.i1(intermediate_wire_3[335]),.i2(intermediate_wire_3[334]),.o(intermediate_reg_3[167])); 
xor_module xor_module_inst_3_32(.clk(clk),.reset(reset),.i1(intermediate_wire_3[333]),.i2(intermediate_wire_3[332]),.o(intermediate_reg_3[166])); 
fsm fsm_inst_3_33(.clk(clk),.reset(reset),.i1(intermediate_wire_3[331]),.i2(intermediate_wire_3[330]),.o(intermediate_reg_3[165])); 
xor_module xor_module_inst_3_34(.clk(clk),.reset(reset),.i1(intermediate_wire_3[329]),.i2(intermediate_wire_3[328]),.o(intermediate_reg_3[164])); 
xor_module xor_module_inst_3_35(.clk(clk),.reset(reset),.i1(intermediate_wire_3[327]),.i2(intermediate_wire_3[326]),.o(intermediate_reg_3[163])); 
xor_module xor_module_inst_3_36(.clk(clk),.reset(reset),.i1(intermediate_wire_3[325]),.i2(intermediate_wire_3[324]),.o(intermediate_reg_3[162])); 
xor_module xor_module_inst_3_37(.clk(clk),.reset(reset),.i1(intermediate_wire_3[323]),.i2(intermediate_wire_3[322]),.o(intermediate_reg_3[161])); 
fsm fsm_inst_3_38(.clk(clk),.reset(reset),.i1(intermediate_wire_3[321]),.i2(intermediate_wire_3[320]),.o(intermediate_reg_3[160])); 
xor_module xor_module_inst_3_39(.clk(clk),.reset(reset),.i1(intermediate_wire_3[319]),.i2(intermediate_wire_3[318]),.o(intermediate_reg_3[159])); 
xor_module xor_module_inst_3_40(.clk(clk),.reset(reset),.i1(intermediate_wire_3[317]),.i2(intermediate_wire_3[316]),.o(intermediate_reg_3[158])); 
fsm fsm_inst_3_41(.clk(clk),.reset(reset),.i1(intermediate_wire_3[315]),.i2(intermediate_wire_3[314]),.o(intermediate_reg_3[157])); 
xor_module xor_module_inst_3_42(.clk(clk),.reset(reset),.i1(intermediate_wire_3[313]),.i2(intermediate_wire_3[312]),.o(intermediate_reg_3[156])); 
xor_module xor_module_inst_3_43(.clk(clk),.reset(reset),.i1(intermediate_wire_3[311]),.i2(intermediate_wire_3[310]),.o(intermediate_reg_3[155])); 
fsm fsm_inst_3_44(.clk(clk),.reset(reset),.i1(intermediate_wire_3[309]),.i2(intermediate_wire_3[308]),.o(intermediate_reg_3[154])); 
fsm fsm_inst_3_45(.clk(clk),.reset(reset),.i1(intermediate_wire_3[307]),.i2(intermediate_wire_3[306]),.o(intermediate_reg_3[153])); 
fsm fsm_inst_3_46(.clk(clk),.reset(reset),.i1(intermediate_wire_3[305]),.i2(intermediate_wire_3[304]),.o(intermediate_reg_3[152])); 
xor_module xor_module_inst_3_47(.clk(clk),.reset(reset),.i1(intermediate_wire_3[303]),.i2(intermediate_wire_3[302]),.o(intermediate_reg_3[151])); 
fsm fsm_inst_3_48(.clk(clk),.reset(reset),.i1(intermediate_wire_3[301]),.i2(intermediate_wire_3[300]),.o(intermediate_reg_3[150])); 
xor_module xor_module_inst_3_49(.clk(clk),.reset(reset),.i1(intermediate_wire_3[299]),.i2(intermediate_wire_3[298]),.o(intermediate_reg_3[149])); 
xor_module xor_module_inst_3_50(.clk(clk),.reset(reset),.i1(intermediate_wire_3[297]),.i2(intermediate_wire_3[296]),.o(intermediate_reg_3[148])); 
xor_module xor_module_inst_3_51(.clk(clk),.reset(reset),.i1(intermediate_wire_3[295]),.i2(intermediate_wire_3[294]),.o(intermediate_reg_3[147])); 
xor_module xor_module_inst_3_52(.clk(clk),.reset(reset),.i1(intermediate_wire_3[293]),.i2(intermediate_wire_3[292]),.o(intermediate_reg_3[146])); 
fsm fsm_inst_3_53(.clk(clk),.reset(reset),.i1(intermediate_wire_3[291]),.i2(intermediate_wire_3[290]),.o(intermediate_reg_3[145])); 
xor_module xor_module_inst_3_54(.clk(clk),.reset(reset),.i1(intermediate_wire_3[289]),.i2(intermediate_wire_3[288]),.o(intermediate_reg_3[144])); 
fsm fsm_inst_3_55(.clk(clk),.reset(reset),.i1(intermediate_wire_3[287]),.i2(intermediate_wire_3[286]),.o(intermediate_reg_3[143])); 
fsm fsm_inst_3_56(.clk(clk),.reset(reset),.i1(intermediate_wire_3[285]),.i2(intermediate_wire_3[284]),.o(intermediate_reg_3[142])); 
fsm fsm_inst_3_57(.clk(clk),.reset(reset),.i1(intermediate_wire_3[283]),.i2(intermediate_wire_3[282]),.o(intermediate_reg_3[141])); 
xor_module xor_module_inst_3_58(.clk(clk),.reset(reset),.i1(intermediate_wire_3[281]),.i2(intermediate_wire_3[280]),.o(intermediate_reg_3[140])); 
xor_module xor_module_inst_3_59(.clk(clk),.reset(reset),.i1(intermediate_wire_3[279]),.i2(intermediate_wire_3[278]),.o(intermediate_reg_3[139])); 
xor_module xor_module_inst_3_60(.clk(clk),.reset(reset),.i1(intermediate_wire_3[277]),.i2(intermediate_wire_3[276]),.o(intermediate_reg_3[138])); 
xor_module xor_module_inst_3_61(.clk(clk),.reset(reset),.i1(intermediate_wire_3[275]),.i2(intermediate_wire_3[274]),.o(intermediate_reg_3[137])); 
fsm fsm_inst_3_62(.clk(clk),.reset(reset),.i1(intermediate_wire_3[273]),.i2(intermediate_wire_3[272]),.o(intermediate_reg_3[136])); 
xor_module xor_module_inst_3_63(.clk(clk),.reset(reset),.i1(intermediate_wire_3[271]),.i2(intermediate_wire_3[270]),.o(intermediate_reg_3[135])); 
fsm fsm_inst_3_64(.clk(clk),.reset(reset),.i1(intermediate_wire_3[269]),.i2(intermediate_wire_3[268]),.o(intermediate_reg_3[134])); 
xor_module xor_module_inst_3_65(.clk(clk),.reset(reset),.i1(intermediate_wire_3[267]),.i2(intermediate_wire_3[266]),.o(intermediate_reg_3[133])); 
xor_module xor_module_inst_3_66(.clk(clk),.reset(reset),.i1(intermediate_wire_3[265]),.i2(intermediate_wire_3[264]),.o(intermediate_reg_3[132])); 
xor_module xor_module_inst_3_67(.clk(clk),.reset(reset),.i1(intermediate_wire_3[263]),.i2(intermediate_wire_3[262]),.o(intermediate_reg_3[131])); 
fsm fsm_inst_3_68(.clk(clk),.reset(reset),.i1(intermediate_wire_3[261]),.i2(intermediate_wire_3[260]),.o(intermediate_reg_3[130])); 
fsm fsm_inst_3_69(.clk(clk),.reset(reset),.i1(intermediate_wire_3[259]),.i2(intermediate_wire_3[258]),.o(intermediate_reg_3[129])); 
xor_module xor_module_inst_3_70(.clk(clk),.reset(reset),.i1(intermediate_wire_3[257]),.i2(intermediate_wire_3[256]),.o(intermediate_reg_3[128])); 
xor_module xor_module_inst_3_71(.clk(clk),.reset(reset),.i1(intermediate_wire_3[255]),.i2(intermediate_wire_3[254]),.o(intermediate_reg_3[127])); 
fsm fsm_inst_3_72(.clk(clk),.reset(reset),.i1(intermediate_wire_3[253]),.i2(intermediate_wire_3[252]),.o(intermediate_reg_3[126])); 
fsm fsm_inst_3_73(.clk(clk),.reset(reset),.i1(intermediate_wire_3[251]),.i2(intermediate_wire_3[250]),.o(intermediate_reg_3[125])); 
fsm fsm_inst_3_74(.clk(clk),.reset(reset),.i1(intermediate_wire_3[249]),.i2(intermediate_wire_3[248]),.o(intermediate_reg_3[124])); 
fsm fsm_inst_3_75(.clk(clk),.reset(reset),.i1(intermediate_wire_3[247]),.i2(intermediate_wire_3[246]),.o(intermediate_reg_3[123])); 
xor_module xor_module_inst_3_76(.clk(clk),.reset(reset),.i1(intermediate_wire_3[245]),.i2(intermediate_wire_3[244]),.o(intermediate_reg_3[122])); 
xor_module xor_module_inst_3_77(.clk(clk),.reset(reset),.i1(intermediate_wire_3[243]),.i2(intermediate_wire_3[242]),.o(intermediate_reg_3[121])); 
xor_module xor_module_inst_3_78(.clk(clk),.reset(reset),.i1(intermediate_wire_3[241]),.i2(intermediate_wire_3[240]),.o(intermediate_reg_3[120])); 
xor_module xor_module_inst_3_79(.clk(clk),.reset(reset),.i1(intermediate_wire_3[239]),.i2(intermediate_wire_3[238]),.o(intermediate_reg_3[119])); 
xor_module xor_module_inst_3_80(.clk(clk),.reset(reset),.i1(intermediate_wire_3[237]),.i2(intermediate_wire_3[236]),.o(intermediate_reg_3[118])); 
xor_module xor_module_inst_3_81(.clk(clk),.reset(reset),.i1(intermediate_wire_3[235]),.i2(intermediate_wire_3[234]),.o(intermediate_reg_3[117])); 
fsm fsm_inst_3_82(.clk(clk),.reset(reset),.i1(intermediate_wire_3[233]),.i2(intermediate_wire_3[232]),.o(intermediate_reg_3[116])); 
fsm fsm_inst_3_83(.clk(clk),.reset(reset),.i1(intermediate_wire_3[231]),.i2(intermediate_wire_3[230]),.o(intermediate_reg_3[115])); 
xor_module xor_module_inst_3_84(.clk(clk),.reset(reset),.i1(intermediate_wire_3[229]),.i2(intermediate_wire_3[228]),.o(intermediate_reg_3[114])); 
xor_module xor_module_inst_3_85(.clk(clk),.reset(reset),.i1(intermediate_wire_3[227]),.i2(intermediate_wire_3[226]),.o(intermediate_reg_3[113])); 
xor_module xor_module_inst_3_86(.clk(clk),.reset(reset),.i1(intermediate_wire_3[225]),.i2(intermediate_wire_3[224]),.o(intermediate_reg_3[112])); 
fsm fsm_inst_3_87(.clk(clk),.reset(reset),.i1(intermediate_wire_3[223]),.i2(intermediate_wire_3[222]),.o(intermediate_reg_3[111])); 
fsm fsm_inst_3_88(.clk(clk),.reset(reset),.i1(intermediate_wire_3[221]),.i2(intermediate_wire_3[220]),.o(intermediate_reg_3[110])); 
xor_module xor_module_inst_3_89(.clk(clk),.reset(reset),.i1(intermediate_wire_3[219]),.i2(intermediate_wire_3[218]),.o(intermediate_reg_3[109])); 
fsm fsm_inst_3_90(.clk(clk),.reset(reset),.i1(intermediate_wire_3[217]),.i2(intermediate_wire_3[216]),.o(intermediate_reg_3[108])); 
fsm fsm_inst_3_91(.clk(clk),.reset(reset),.i1(intermediate_wire_3[215]),.i2(intermediate_wire_3[214]),.o(intermediate_reg_3[107])); 
xor_module xor_module_inst_3_92(.clk(clk),.reset(reset),.i1(intermediate_wire_3[213]),.i2(intermediate_wire_3[212]),.o(intermediate_reg_3[106])); 
fsm fsm_inst_3_93(.clk(clk),.reset(reset),.i1(intermediate_wire_3[211]),.i2(intermediate_wire_3[210]),.o(intermediate_reg_3[105])); 
fsm fsm_inst_3_94(.clk(clk),.reset(reset),.i1(intermediate_wire_3[209]),.i2(intermediate_wire_3[208]),.o(intermediate_reg_3[104])); 
xor_module xor_module_inst_3_95(.clk(clk),.reset(reset),.i1(intermediate_wire_3[207]),.i2(intermediate_wire_3[206]),.o(intermediate_reg_3[103])); 
xor_module xor_module_inst_3_96(.clk(clk),.reset(reset),.i1(intermediate_wire_3[205]),.i2(intermediate_wire_3[204]),.o(intermediate_reg_3[102])); 
fsm fsm_inst_3_97(.clk(clk),.reset(reset),.i1(intermediate_wire_3[203]),.i2(intermediate_wire_3[202]),.o(intermediate_reg_3[101])); 
fsm fsm_inst_3_98(.clk(clk),.reset(reset),.i1(intermediate_wire_3[201]),.i2(intermediate_wire_3[200]),.o(intermediate_reg_3[100])); 
fsm fsm_inst_3_99(.clk(clk),.reset(reset),.i1(intermediate_wire_3[199]),.i2(intermediate_wire_3[198]),.o(intermediate_reg_3[99])); 
fsm fsm_inst_3_100(.clk(clk),.reset(reset),.i1(intermediate_wire_3[197]),.i2(intermediate_wire_3[196]),.o(intermediate_reg_3[98])); 
xor_module xor_module_inst_3_101(.clk(clk),.reset(reset),.i1(intermediate_wire_3[195]),.i2(intermediate_wire_3[194]),.o(intermediate_reg_3[97])); 
fsm fsm_inst_3_102(.clk(clk),.reset(reset),.i1(intermediate_wire_3[193]),.i2(intermediate_wire_3[192]),.o(intermediate_reg_3[96])); 
xor_module xor_module_inst_3_103(.clk(clk),.reset(reset),.i1(intermediate_wire_3[191]),.i2(intermediate_wire_3[190]),.o(intermediate_reg_3[95])); 
fsm fsm_inst_3_104(.clk(clk),.reset(reset),.i1(intermediate_wire_3[189]),.i2(intermediate_wire_3[188]),.o(intermediate_reg_3[94])); 
fsm fsm_inst_3_105(.clk(clk),.reset(reset),.i1(intermediate_wire_3[187]),.i2(intermediate_wire_3[186]),.o(intermediate_reg_3[93])); 
xor_module xor_module_inst_3_106(.clk(clk),.reset(reset),.i1(intermediate_wire_3[185]),.i2(intermediate_wire_3[184]),.o(intermediate_reg_3[92])); 
fsm fsm_inst_3_107(.clk(clk),.reset(reset),.i1(intermediate_wire_3[183]),.i2(intermediate_wire_3[182]),.o(intermediate_reg_3[91])); 
fsm fsm_inst_3_108(.clk(clk),.reset(reset),.i1(intermediate_wire_3[181]),.i2(intermediate_wire_3[180]),.o(intermediate_reg_3[90])); 
xor_module xor_module_inst_3_109(.clk(clk),.reset(reset),.i1(intermediate_wire_3[179]),.i2(intermediate_wire_3[178]),.o(intermediate_reg_3[89])); 
xor_module xor_module_inst_3_110(.clk(clk),.reset(reset),.i1(intermediate_wire_3[177]),.i2(intermediate_wire_3[176]),.o(intermediate_reg_3[88])); 
fsm fsm_inst_3_111(.clk(clk),.reset(reset),.i1(intermediate_wire_3[175]),.i2(intermediate_wire_3[174]),.o(intermediate_reg_3[87])); 
xor_module xor_module_inst_3_112(.clk(clk),.reset(reset),.i1(intermediate_wire_3[173]),.i2(intermediate_wire_3[172]),.o(intermediate_reg_3[86])); 
xor_module xor_module_inst_3_113(.clk(clk),.reset(reset),.i1(intermediate_wire_3[171]),.i2(intermediate_wire_3[170]),.o(intermediate_reg_3[85])); 
xor_module xor_module_inst_3_114(.clk(clk),.reset(reset),.i1(intermediate_wire_3[169]),.i2(intermediate_wire_3[168]),.o(intermediate_reg_3[84])); 
fsm fsm_inst_3_115(.clk(clk),.reset(reset),.i1(intermediate_wire_3[167]),.i2(intermediate_wire_3[166]),.o(intermediate_reg_3[83])); 
xor_module xor_module_inst_3_116(.clk(clk),.reset(reset),.i1(intermediate_wire_3[165]),.i2(intermediate_wire_3[164]),.o(intermediate_reg_3[82])); 
fsm fsm_inst_3_117(.clk(clk),.reset(reset),.i1(intermediate_wire_3[163]),.i2(intermediate_wire_3[162]),.o(intermediate_reg_3[81])); 
fsm fsm_inst_3_118(.clk(clk),.reset(reset),.i1(intermediate_wire_3[161]),.i2(intermediate_wire_3[160]),.o(intermediate_reg_3[80])); 
fsm fsm_inst_3_119(.clk(clk),.reset(reset),.i1(intermediate_wire_3[159]),.i2(intermediate_wire_3[158]),.o(intermediate_reg_3[79])); 
fsm fsm_inst_3_120(.clk(clk),.reset(reset),.i1(intermediate_wire_3[157]),.i2(intermediate_wire_3[156]),.o(intermediate_reg_3[78])); 
xor_module xor_module_inst_3_121(.clk(clk),.reset(reset),.i1(intermediate_wire_3[155]),.i2(intermediate_wire_3[154]),.o(intermediate_reg_3[77])); 
xor_module xor_module_inst_3_122(.clk(clk),.reset(reset),.i1(intermediate_wire_3[153]),.i2(intermediate_wire_3[152]),.o(intermediate_reg_3[76])); 
fsm fsm_inst_3_123(.clk(clk),.reset(reset),.i1(intermediate_wire_3[151]),.i2(intermediate_wire_3[150]),.o(intermediate_reg_3[75])); 
xor_module xor_module_inst_3_124(.clk(clk),.reset(reset),.i1(intermediate_wire_3[149]),.i2(intermediate_wire_3[148]),.o(intermediate_reg_3[74])); 
fsm fsm_inst_3_125(.clk(clk),.reset(reset),.i1(intermediate_wire_3[147]),.i2(intermediate_wire_3[146]),.o(intermediate_reg_3[73])); 
fsm fsm_inst_3_126(.clk(clk),.reset(reset),.i1(intermediate_wire_3[145]),.i2(intermediate_wire_3[144]),.o(intermediate_reg_3[72])); 
fsm fsm_inst_3_127(.clk(clk),.reset(reset),.i1(intermediate_wire_3[143]),.i2(intermediate_wire_3[142]),.o(intermediate_reg_3[71])); 
fsm fsm_inst_3_128(.clk(clk),.reset(reset),.i1(intermediate_wire_3[141]),.i2(intermediate_wire_3[140]),.o(intermediate_reg_3[70])); 
xor_module xor_module_inst_3_129(.clk(clk),.reset(reset),.i1(intermediate_wire_3[139]),.i2(intermediate_wire_3[138]),.o(intermediate_reg_3[69])); 
fsm fsm_inst_3_130(.clk(clk),.reset(reset),.i1(intermediate_wire_3[137]),.i2(intermediate_wire_3[136]),.o(intermediate_reg_3[68])); 
fsm fsm_inst_3_131(.clk(clk),.reset(reset),.i1(intermediate_wire_3[135]),.i2(intermediate_wire_3[134]),.o(intermediate_reg_3[67])); 
fsm fsm_inst_3_132(.clk(clk),.reset(reset),.i1(intermediate_wire_3[133]),.i2(intermediate_wire_3[132]),.o(intermediate_reg_3[66])); 
fsm fsm_inst_3_133(.clk(clk),.reset(reset),.i1(intermediate_wire_3[131]),.i2(intermediate_wire_3[130]),.o(intermediate_reg_3[65])); 
xor_module xor_module_inst_3_134(.clk(clk),.reset(reset),.i1(intermediate_wire_3[129]),.i2(intermediate_wire_3[128]),.o(intermediate_reg_3[64])); 
fsm fsm_inst_3_135(.clk(clk),.reset(reset),.i1(intermediate_wire_3[127]),.i2(intermediate_wire_3[126]),.o(intermediate_reg_3[63])); 
fsm fsm_inst_3_136(.clk(clk),.reset(reset),.i1(intermediate_wire_3[125]),.i2(intermediate_wire_3[124]),.o(intermediate_reg_3[62])); 
xor_module xor_module_inst_3_137(.clk(clk),.reset(reset),.i1(intermediate_wire_3[123]),.i2(intermediate_wire_3[122]),.o(intermediate_reg_3[61])); 
fsm fsm_inst_3_138(.clk(clk),.reset(reset),.i1(intermediate_wire_3[121]),.i2(intermediate_wire_3[120]),.o(intermediate_reg_3[60])); 
xor_module xor_module_inst_3_139(.clk(clk),.reset(reset),.i1(intermediate_wire_3[119]),.i2(intermediate_wire_3[118]),.o(intermediate_reg_3[59])); 
fsm fsm_inst_3_140(.clk(clk),.reset(reset),.i1(intermediate_wire_3[117]),.i2(intermediate_wire_3[116]),.o(intermediate_reg_3[58])); 
xor_module xor_module_inst_3_141(.clk(clk),.reset(reset),.i1(intermediate_wire_3[115]),.i2(intermediate_wire_3[114]),.o(intermediate_reg_3[57])); 
fsm fsm_inst_3_142(.clk(clk),.reset(reset),.i1(intermediate_wire_3[113]),.i2(intermediate_wire_3[112]),.o(intermediate_reg_3[56])); 
fsm fsm_inst_3_143(.clk(clk),.reset(reset),.i1(intermediate_wire_3[111]),.i2(intermediate_wire_3[110]),.o(intermediate_reg_3[55])); 
fsm fsm_inst_3_144(.clk(clk),.reset(reset),.i1(intermediate_wire_3[109]),.i2(intermediate_wire_3[108]),.o(intermediate_reg_3[54])); 
xor_module xor_module_inst_3_145(.clk(clk),.reset(reset),.i1(intermediate_wire_3[107]),.i2(intermediate_wire_3[106]),.o(intermediate_reg_3[53])); 
xor_module xor_module_inst_3_146(.clk(clk),.reset(reset),.i1(intermediate_wire_3[105]),.i2(intermediate_wire_3[104]),.o(intermediate_reg_3[52])); 
xor_module xor_module_inst_3_147(.clk(clk),.reset(reset),.i1(intermediate_wire_3[103]),.i2(intermediate_wire_3[102]),.o(intermediate_reg_3[51])); 
xor_module xor_module_inst_3_148(.clk(clk),.reset(reset),.i1(intermediate_wire_3[101]),.i2(intermediate_wire_3[100]),.o(intermediate_reg_3[50])); 
fsm fsm_inst_3_149(.clk(clk),.reset(reset),.i1(intermediate_wire_3[99]),.i2(intermediate_wire_3[98]),.o(intermediate_reg_3[49])); 
xor_module xor_module_inst_3_150(.clk(clk),.reset(reset),.i1(intermediate_wire_3[97]),.i2(intermediate_wire_3[96]),.o(intermediate_reg_3[48])); 
xor_module xor_module_inst_3_151(.clk(clk),.reset(reset),.i1(intermediate_wire_3[95]),.i2(intermediate_wire_3[94]),.o(intermediate_reg_3[47])); 
fsm fsm_inst_3_152(.clk(clk),.reset(reset),.i1(intermediate_wire_3[93]),.i2(intermediate_wire_3[92]),.o(intermediate_reg_3[46])); 
xor_module xor_module_inst_3_153(.clk(clk),.reset(reset),.i1(intermediate_wire_3[91]),.i2(intermediate_wire_3[90]),.o(intermediate_reg_3[45])); 
fsm fsm_inst_3_154(.clk(clk),.reset(reset),.i1(intermediate_wire_3[89]),.i2(intermediate_wire_3[88]),.o(intermediate_reg_3[44])); 
xor_module xor_module_inst_3_155(.clk(clk),.reset(reset),.i1(intermediate_wire_3[87]),.i2(intermediate_wire_3[86]),.o(intermediate_reg_3[43])); 
xor_module xor_module_inst_3_156(.clk(clk),.reset(reset),.i1(intermediate_wire_3[85]),.i2(intermediate_wire_3[84]),.o(intermediate_reg_3[42])); 
fsm fsm_inst_3_157(.clk(clk),.reset(reset),.i1(intermediate_wire_3[83]),.i2(intermediate_wire_3[82]),.o(intermediate_reg_3[41])); 
fsm fsm_inst_3_158(.clk(clk),.reset(reset),.i1(intermediate_wire_3[81]),.i2(intermediate_wire_3[80]),.o(intermediate_reg_3[40])); 
fsm fsm_inst_3_159(.clk(clk),.reset(reset),.i1(intermediate_wire_3[79]),.i2(intermediate_wire_3[78]),.o(intermediate_reg_3[39])); 
xor_module xor_module_inst_3_160(.clk(clk),.reset(reset),.i1(intermediate_wire_3[77]),.i2(intermediate_wire_3[76]),.o(intermediate_reg_3[38])); 
fsm fsm_inst_3_161(.clk(clk),.reset(reset),.i1(intermediate_wire_3[75]),.i2(intermediate_wire_3[74]),.o(intermediate_reg_3[37])); 
xor_module xor_module_inst_3_162(.clk(clk),.reset(reset),.i1(intermediate_wire_3[73]),.i2(intermediate_wire_3[72]),.o(intermediate_reg_3[36])); 
fsm fsm_inst_3_163(.clk(clk),.reset(reset),.i1(intermediate_wire_3[71]),.i2(intermediate_wire_3[70]),.o(intermediate_reg_3[35])); 
fsm fsm_inst_3_164(.clk(clk),.reset(reset),.i1(intermediate_wire_3[69]),.i2(intermediate_wire_3[68]),.o(intermediate_reg_3[34])); 
xor_module xor_module_inst_3_165(.clk(clk),.reset(reset),.i1(intermediate_wire_3[67]),.i2(intermediate_wire_3[66]),.o(intermediate_reg_3[33])); 
xor_module xor_module_inst_3_166(.clk(clk),.reset(reset),.i1(intermediate_wire_3[65]),.i2(intermediate_wire_3[64]),.o(intermediate_reg_3[32])); 
fsm fsm_inst_3_167(.clk(clk),.reset(reset),.i1(intermediate_wire_3[63]),.i2(intermediate_wire_3[62]),.o(intermediate_reg_3[31])); 
xor_module xor_module_inst_3_168(.clk(clk),.reset(reset),.i1(intermediate_wire_3[61]),.i2(intermediate_wire_3[60]),.o(intermediate_reg_3[30])); 
fsm fsm_inst_3_169(.clk(clk),.reset(reset),.i1(intermediate_wire_3[59]),.i2(intermediate_wire_3[58]),.o(intermediate_reg_3[29])); 
xor_module xor_module_inst_3_170(.clk(clk),.reset(reset),.i1(intermediate_wire_3[57]),.i2(intermediate_wire_3[56]),.o(intermediate_reg_3[28])); 
fsm fsm_inst_3_171(.clk(clk),.reset(reset),.i1(intermediate_wire_3[55]),.i2(intermediate_wire_3[54]),.o(intermediate_reg_3[27])); 
xor_module xor_module_inst_3_172(.clk(clk),.reset(reset),.i1(intermediate_wire_3[53]),.i2(intermediate_wire_3[52]),.o(intermediate_reg_3[26])); 
xor_module xor_module_inst_3_173(.clk(clk),.reset(reset),.i1(intermediate_wire_3[51]),.i2(intermediate_wire_3[50]),.o(intermediate_reg_3[25])); 
fsm fsm_inst_3_174(.clk(clk),.reset(reset),.i1(intermediate_wire_3[49]),.i2(intermediate_wire_3[48]),.o(intermediate_reg_3[24])); 
fsm fsm_inst_3_175(.clk(clk),.reset(reset),.i1(intermediate_wire_3[47]),.i2(intermediate_wire_3[46]),.o(intermediate_reg_3[23])); 
xor_module xor_module_inst_3_176(.clk(clk),.reset(reset),.i1(intermediate_wire_3[45]),.i2(intermediate_wire_3[44]),.o(intermediate_reg_3[22])); 
fsm fsm_inst_3_177(.clk(clk),.reset(reset),.i1(intermediate_wire_3[43]),.i2(intermediate_wire_3[42]),.o(intermediate_reg_3[21])); 
fsm fsm_inst_3_178(.clk(clk),.reset(reset),.i1(intermediate_wire_3[41]),.i2(intermediate_wire_3[40]),.o(intermediate_reg_3[20])); 
fsm fsm_inst_3_179(.clk(clk),.reset(reset),.i1(intermediate_wire_3[39]),.i2(intermediate_wire_3[38]),.o(intermediate_reg_3[19])); 
xor_module xor_module_inst_3_180(.clk(clk),.reset(reset),.i1(intermediate_wire_3[37]),.i2(intermediate_wire_3[36]),.o(intermediate_reg_3[18])); 
fsm fsm_inst_3_181(.clk(clk),.reset(reset),.i1(intermediate_wire_3[35]),.i2(intermediate_wire_3[34]),.o(intermediate_reg_3[17])); 
xor_module xor_module_inst_3_182(.clk(clk),.reset(reset),.i1(intermediate_wire_3[33]),.i2(intermediate_wire_3[32]),.o(intermediate_reg_3[16])); 
xor_module xor_module_inst_3_183(.clk(clk),.reset(reset),.i1(intermediate_wire_3[31]),.i2(intermediate_wire_3[30]),.o(intermediate_reg_3[15])); 
xor_module xor_module_inst_3_184(.clk(clk),.reset(reset),.i1(intermediate_wire_3[29]),.i2(intermediate_wire_3[28]),.o(intermediate_reg_3[14])); 
fsm fsm_inst_3_185(.clk(clk),.reset(reset),.i1(intermediate_wire_3[27]),.i2(intermediate_wire_3[26]),.o(intermediate_reg_3[13])); 
fsm fsm_inst_3_186(.clk(clk),.reset(reset),.i1(intermediate_wire_3[25]),.i2(intermediate_wire_3[24]),.o(intermediate_reg_3[12])); 
fsm fsm_inst_3_187(.clk(clk),.reset(reset),.i1(intermediate_wire_3[23]),.i2(intermediate_wire_3[22]),.o(intermediate_reg_3[11])); 
xor_module xor_module_inst_3_188(.clk(clk),.reset(reset),.i1(intermediate_wire_3[21]),.i2(intermediate_wire_3[20]),.o(intermediate_reg_3[10])); 
fsm fsm_inst_3_189(.clk(clk),.reset(reset),.i1(intermediate_wire_3[19]),.i2(intermediate_wire_3[18]),.o(intermediate_reg_3[9])); 
fsm fsm_inst_3_190(.clk(clk),.reset(reset),.i1(intermediate_wire_3[17]),.i2(intermediate_wire_3[16]),.o(intermediate_reg_3[8])); 
fsm fsm_inst_3_191(.clk(clk),.reset(reset),.i1(intermediate_wire_3[15]),.i2(intermediate_wire_3[14]),.o(intermediate_reg_3[7])); 
fsm fsm_inst_3_192(.clk(clk),.reset(reset),.i1(intermediate_wire_3[13]),.i2(intermediate_wire_3[12]),.o(intermediate_reg_3[6])); 
xor_module xor_module_inst_3_193(.clk(clk),.reset(reset),.i1(intermediate_wire_3[11]),.i2(intermediate_wire_3[10]),.o(intermediate_reg_3[5])); 
xor_module xor_module_inst_3_194(.clk(clk),.reset(reset),.i1(intermediate_wire_3[9]),.i2(intermediate_wire_3[8]),.o(intermediate_reg_3[4])); 
xor_module xor_module_inst_3_195(.clk(clk),.reset(reset),.i1(intermediate_wire_3[7]),.i2(intermediate_wire_3[6]),.o(intermediate_reg_3[3])); 
xor_module xor_module_inst_3_196(.clk(clk),.reset(reset),.i1(intermediate_wire_3[5]),.i2(intermediate_wire_3[4]),.o(intermediate_reg_3[2])); 
xor_module xor_module_inst_3_197(.clk(clk),.reset(reset),.i1(intermediate_wire_3[3]),.i2(intermediate_wire_3[2]),.o(intermediate_reg_3[1])); 
fsm fsm_inst_3_198(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1]),.i2(intermediate_wire_3[0]),.o(intermediate_reg_3[0])); 
wire [197:0]intermediate_wire_4; 
assign intermediate_wire_4[197] = intermediate_reg_3[198]^intermediate_reg_3[197] ; 
assign intermediate_wire_4[196:0] = intermediate_reg_3[196:0] ; 
reg [98:0]intermediate_reg_4; 
 
fsm fsm_inst_4_0(.clk(clk),.reset(reset),.i1(intermediate_wire_4[197]),.i2(intermediate_wire_4[196]),.o(intermediate_reg_4[98])); 
fsm fsm_inst_4_1(.clk(clk),.reset(reset),.i1(intermediate_wire_4[195]),.i2(intermediate_wire_4[194]),.o(intermediate_reg_4[97])); 
fsm fsm_inst_4_2(.clk(clk),.reset(reset),.i1(intermediate_wire_4[193]),.i2(intermediate_wire_4[192]),.o(intermediate_reg_4[96])); 
xor_module xor_module_inst_4_3(.clk(clk),.reset(reset),.i1(intermediate_wire_4[191]),.i2(intermediate_wire_4[190]),.o(intermediate_reg_4[95])); 
xor_module xor_module_inst_4_4(.clk(clk),.reset(reset),.i1(intermediate_wire_4[189]),.i2(intermediate_wire_4[188]),.o(intermediate_reg_4[94])); 
fsm fsm_inst_4_5(.clk(clk),.reset(reset),.i1(intermediate_wire_4[187]),.i2(intermediate_wire_4[186]),.o(intermediate_reg_4[93])); 
xor_module xor_module_inst_4_6(.clk(clk),.reset(reset),.i1(intermediate_wire_4[185]),.i2(intermediate_wire_4[184]),.o(intermediate_reg_4[92])); 
xor_module xor_module_inst_4_7(.clk(clk),.reset(reset),.i1(intermediate_wire_4[183]),.i2(intermediate_wire_4[182]),.o(intermediate_reg_4[91])); 
xor_module xor_module_inst_4_8(.clk(clk),.reset(reset),.i1(intermediate_wire_4[181]),.i2(intermediate_wire_4[180]),.o(intermediate_reg_4[90])); 
fsm fsm_inst_4_9(.clk(clk),.reset(reset),.i1(intermediate_wire_4[179]),.i2(intermediate_wire_4[178]),.o(intermediate_reg_4[89])); 
xor_module xor_module_inst_4_10(.clk(clk),.reset(reset),.i1(intermediate_wire_4[177]),.i2(intermediate_wire_4[176]),.o(intermediate_reg_4[88])); 
xor_module xor_module_inst_4_11(.clk(clk),.reset(reset),.i1(intermediate_wire_4[175]),.i2(intermediate_wire_4[174]),.o(intermediate_reg_4[87])); 
xor_module xor_module_inst_4_12(.clk(clk),.reset(reset),.i1(intermediate_wire_4[173]),.i2(intermediate_wire_4[172]),.o(intermediate_reg_4[86])); 
fsm fsm_inst_4_13(.clk(clk),.reset(reset),.i1(intermediate_wire_4[171]),.i2(intermediate_wire_4[170]),.o(intermediate_reg_4[85])); 
xor_module xor_module_inst_4_14(.clk(clk),.reset(reset),.i1(intermediate_wire_4[169]),.i2(intermediate_wire_4[168]),.o(intermediate_reg_4[84])); 
fsm fsm_inst_4_15(.clk(clk),.reset(reset),.i1(intermediate_wire_4[167]),.i2(intermediate_wire_4[166]),.o(intermediate_reg_4[83])); 
fsm fsm_inst_4_16(.clk(clk),.reset(reset),.i1(intermediate_wire_4[165]),.i2(intermediate_wire_4[164]),.o(intermediate_reg_4[82])); 
fsm fsm_inst_4_17(.clk(clk),.reset(reset),.i1(intermediate_wire_4[163]),.i2(intermediate_wire_4[162]),.o(intermediate_reg_4[81])); 
fsm fsm_inst_4_18(.clk(clk),.reset(reset),.i1(intermediate_wire_4[161]),.i2(intermediate_wire_4[160]),.o(intermediate_reg_4[80])); 
xor_module xor_module_inst_4_19(.clk(clk),.reset(reset),.i1(intermediate_wire_4[159]),.i2(intermediate_wire_4[158]),.o(intermediate_reg_4[79])); 
xor_module xor_module_inst_4_20(.clk(clk),.reset(reset),.i1(intermediate_wire_4[157]),.i2(intermediate_wire_4[156]),.o(intermediate_reg_4[78])); 
xor_module xor_module_inst_4_21(.clk(clk),.reset(reset),.i1(intermediate_wire_4[155]),.i2(intermediate_wire_4[154]),.o(intermediate_reg_4[77])); 
xor_module xor_module_inst_4_22(.clk(clk),.reset(reset),.i1(intermediate_wire_4[153]),.i2(intermediate_wire_4[152]),.o(intermediate_reg_4[76])); 
xor_module xor_module_inst_4_23(.clk(clk),.reset(reset),.i1(intermediate_wire_4[151]),.i2(intermediate_wire_4[150]),.o(intermediate_reg_4[75])); 
fsm fsm_inst_4_24(.clk(clk),.reset(reset),.i1(intermediate_wire_4[149]),.i2(intermediate_wire_4[148]),.o(intermediate_reg_4[74])); 
xor_module xor_module_inst_4_25(.clk(clk),.reset(reset),.i1(intermediate_wire_4[147]),.i2(intermediate_wire_4[146]),.o(intermediate_reg_4[73])); 
fsm fsm_inst_4_26(.clk(clk),.reset(reset),.i1(intermediate_wire_4[145]),.i2(intermediate_wire_4[144]),.o(intermediate_reg_4[72])); 
xor_module xor_module_inst_4_27(.clk(clk),.reset(reset),.i1(intermediate_wire_4[143]),.i2(intermediate_wire_4[142]),.o(intermediate_reg_4[71])); 
xor_module xor_module_inst_4_28(.clk(clk),.reset(reset),.i1(intermediate_wire_4[141]),.i2(intermediate_wire_4[140]),.o(intermediate_reg_4[70])); 
fsm fsm_inst_4_29(.clk(clk),.reset(reset),.i1(intermediate_wire_4[139]),.i2(intermediate_wire_4[138]),.o(intermediate_reg_4[69])); 
fsm fsm_inst_4_30(.clk(clk),.reset(reset),.i1(intermediate_wire_4[137]),.i2(intermediate_wire_4[136]),.o(intermediate_reg_4[68])); 
fsm fsm_inst_4_31(.clk(clk),.reset(reset),.i1(intermediate_wire_4[135]),.i2(intermediate_wire_4[134]),.o(intermediate_reg_4[67])); 
xor_module xor_module_inst_4_32(.clk(clk),.reset(reset),.i1(intermediate_wire_4[133]),.i2(intermediate_wire_4[132]),.o(intermediate_reg_4[66])); 
xor_module xor_module_inst_4_33(.clk(clk),.reset(reset),.i1(intermediate_wire_4[131]),.i2(intermediate_wire_4[130]),.o(intermediate_reg_4[65])); 
xor_module xor_module_inst_4_34(.clk(clk),.reset(reset),.i1(intermediate_wire_4[129]),.i2(intermediate_wire_4[128]),.o(intermediate_reg_4[64])); 
fsm fsm_inst_4_35(.clk(clk),.reset(reset),.i1(intermediate_wire_4[127]),.i2(intermediate_wire_4[126]),.o(intermediate_reg_4[63])); 
fsm fsm_inst_4_36(.clk(clk),.reset(reset),.i1(intermediate_wire_4[125]),.i2(intermediate_wire_4[124]),.o(intermediate_reg_4[62])); 
xor_module xor_module_inst_4_37(.clk(clk),.reset(reset),.i1(intermediate_wire_4[123]),.i2(intermediate_wire_4[122]),.o(intermediate_reg_4[61])); 
xor_module xor_module_inst_4_38(.clk(clk),.reset(reset),.i1(intermediate_wire_4[121]),.i2(intermediate_wire_4[120]),.o(intermediate_reg_4[60])); 
fsm fsm_inst_4_39(.clk(clk),.reset(reset),.i1(intermediate_wire_4[119]),.i2(intermediate_wire_4[118]),.o(intermediate_reg_4[59])); 
fsm fsm_inst_4_40(.clk(clk),.reset(reset),.i1(intermediate_wire_4[117]),.i2(intermediate_wire_4[116]),.o(intermediate_reg_4[58])); 
fsm fsm_inst_4_41(.clk(clk),.reset(reset),.i1(intermediate_wire_4[115]),.i2(intermediate_wire_4[114]),.o(intermediate_reg_4[57])); 
xor_module xor_module_inst_4_42(.clk(clk),.reset(reset),.i1(intermediate_wire_4[113]),.i2(intermediate_wire_4[112]),.o(intermediate_reg_4[56])); 
xor_module xor_module_inst_4_43(.clk(clk),.reset(reset),.i1(intermediate_wire_4[111]),.i2(intermediate_wire_4[110]),.o(intermediate_reg_4[55])); 
fsm fsm_inst_4_44(.clk(clk),.reset(reset),.i1(intermediate_wire_4[109]),.i2(intermediate_wire_4[108]),.o(intermediate_reg_4[54])); 
fsm fsm_inst_4_45(.clk(clk),.reset(reset),.i1(intermediate_wire_4[107]),.i2(intermediate_wire_4[106]),.o(intermediate_reg_4[53])); 
xor_module xor_module_inst_4_46(.clk(clk),.reset(reset),.i1(intermediate_wire_4[105]),.i2(intermediate_wire_4[104]),.o(intermediate_reg_4[52])); 
fsm fsm_inst_4_47(.clk(clk),.reset(reset),.i1(intermediate_wire_4[103]),.i2(intermediate_wire_4[102]),.o(intermediate_reg_4[51])); 
xor_module xor_module_inst_4_48(.clk(clk),.reset(reset),.i1(intermediate_wire_4[101]),.i2(intermediate_wire_4[100]),.o(intermediate_reg_4[50])); 
xor_module xor_module_inst_4_49(.clk(clk),.reset(reset),.i1(intermediate_wire_4[99]),.i2(intermediate_wire_4[98]),.o(intermediate_reg_4[49])); 
fsm fsm_inst_4_50(.clk(clk),.reset(reset),.i1(intermediate_wire_4[97]),.i2(intermediate_wire_4[96]),.o(intermediate_reg_4[48])); 
xor_module xor_module_inst_4_51(.clk(clk),.reset(reset),.i1(intermediate_wire_4[95]),.i2(intermediate_wire_4[94]),.o(intermediate_reg_4[47])); 
xor_module xor_module_inst_4_52(.clk(clk),.reset(reset),.i1(intermediate_wire_4[93]),.i2(intermediate_wire_4[92]),.o(intermediate_reg_4[46])); 
xor_module xor_module_inst_4_53(.clk(clk),.reset(reset),.i1(intermediate_wire_4[91]),.i2(intermediate_wire_4[90]),.o(intermediate_reg_4[45])); 
xor_module xor_module_inst_4_54(.clk(clk),.reset(reset),.i1(intermediate_wire_4[89]),.i2(intermediate_wire_4[88]),.o(intermediate_reg_4[44])); 
fsm fsm_inst_4_55(.clk(clk),.reset(reset),.i1(intermediate_wire_4[87]),.i2(intermediate_wire_4[86]),.o(intermediate_reg_4[43])); 
fsm fsm_inst_4_56(.clk(clk),.reset(reset),.i1(intermediate_wire_4[85]),.i2(intermediate_wire_4[84]),.o(intermediate_reg_4[42])); 
xor_module xor_module_inst_4_57(.clk(clk),.reset(reset),.i1(intermediate_wire_4[83]),.i2(intermediate_wire_4[82]),.o(intermediate_reg_4[41])); 
fsm fsm_inst_4_58(.clk(clk),.reset(reset),.i1(intermediate_wire_4[81]),.i2(intermediate_wire_4[80]),.o(intermediate_reg_4[40])); 
xor_module xor_module_inst_4_59(.clk(clk),.reset(reset),.i1(intermediate_wire_4[79]),.i2(intermediate_wire_4[78]),.o(intermediate_reg_4[39])); 
fsm fsm_inst_4_60(.clk(clk),.reset(reset),.i1(intermediate_wire_4[77]),.i2(intermediate_wire_4[76]),.o(intermediate_reg_4[38])); 
xor_module xor_module_inst_4_61(.clk(clk),.reset(reset),.i1(intermediate_wire_4[75]),.i2(intermediate_wire_4[74]),.o(intermediate_reg_4[37])); 
xor_module xor_module_inst_4_62(.clk(clk),.reset(reset),.i1(intermediate_wire_4[73]),.i2(intermediate_wire_4[72]),.o(intermediate_reg_4[36])); 
fsm fsm_inst_4_63(.clk(clk),.reset(reset),.i1(intermediate_wire_4[71]),.i2(intermediate_wire_4[70]),.o(intermediate_reg_4[35])); 
xor_module xor_module_inst_4_64(.clk(clk),.reset(reset),.i1(intermediate_wire_4[69]),.i2(intermediate_wire_4[68]),.o(intermediate_reg_4[34])); 
fsm fsm_inst_4_65(.clk(clk),.reset(reset),.i1(intermediate_wire_4[67]),.i2(intermediate_wire_4[66]),.o(intermediate_reg_4[33])); 
fsm fsm_inst_4_66(.clk(clk),.reset(reset),.i1(intermediate_wire_4[65]),.i2(intermediate_wire_4[64]),.o(intermediate_reg_4[32])); 
xor_module xor_module_inst_4_67(.clk(clk),.reset(reset),.i1(intermediate_wire_4[63]),.i2(intermediate_wire_4[62]),.o(intermediate_reg_4[31])); 
xor_module xor_module_inst_4_68(.clk(clk),.reset(reset),.i1(intermediate_wire_4[61]),.i2(intermediate_wire_4[60]),.o(intermediate_reg_4[30])); 
fsm fsm_inst_4_69(.clk(clk),.reset(reset),.i1(intermediate_wire_4[59]),.i2(intermediate_wire_4[58]),.o(intermediate_reg_4[29])); 
xor_module xor_module_inst_4_70(.clk(clk),.reset(reset),.i1(intermediate_wire_4[57]),.i2(intermediate_wire_4[56]),.o(intermediate_reg_4[28])); 
fsm fsm_inst_4_71(.clk(clk),.reset(reset),.i1(intermediate_wire_4[55]),.i2(intermediate_wire_4[54]),.o(intermediate_reg_4[27])); 
fsm fsm_inst_4_72(.clk(clk),.reset(reset),.i1(intermediate_wire_4[53]),.i2(intermediate_wire_4[52]),.o(intermediate_reg_4[26])); 
fsm fsm_inst_4_73(.clk(clk),.reset(reset),.i1(intermediate_wire_4[51]),.i2(intermediate_wire_4[50]),.o(intermediate_reg_4[25])); 
fsm fsm_inst_4_74(.clk(clk),.reset(reset),.i1(intermediate_wire_4[49]),.i2(intermediate_wire_4[48]),.o(intermediate_reg_4[24])); 
xor_module xor_module_inst_4_75(.clk(clk),.reset(reset),.i1(intermediate_wire_4[47]),.i2(intermediate_wire_4[46]),.o(intermediate_reg_4[23])); 
fsm fsm_inst_4_76(.clk(clk),.reset(reset),.i1(intermediate_wire_4[45]),.i2(intermediate_wire_4[44]),.o(intermediate_reg_4[22])); 
fsm fsm_inst_4_77(.clk(clk),.reset(reset),.i1(intermediate_wire_4[43]),.i2(intermediate_wire_4[42]),.o(intermediate_reg_4[21])); 
xor_module xor_module_inst_4_78(.clk(clk),.reset(reset),.i1(intermediate_wire_4[41]),.i2(intermediate_wire_4[40]),.o(intermediate_reg_4[20])); 
xor_module xor_module_inst_4_79(.clk(clk),.reset(reset),.i1(intermediate_wire_4[39]),.i2(intermediate_wire_4[38]),.o(intermediate_reg_4[19])); 
xor_module xor_module_inst_4_80(.clk(clk),.reset(reset),.i1(intermediate_wire_4[37]),.i2(intermediate_wire_4[36]),.o(intermediate_reg_4[18])); 
xor_module xor_module_inst_4_81(.clk(clk),.reset(reset),.i1(intermediate_wire_4[35]),.i2(intermediate_wire_4[34]),.o(intermediate_reg_4[17])); 
xor_module xor_module_inst_4_82(.clk(clk),.reset(reset),.i1(intermediate_wire_4[33]),.i2(intermediate_wire_4[32]),.o(intermediate_reg_4[16])); 
fsm fsm_inst_4_83(.clk(clk),.reset(reset),.i1(intermediate_wire_4[31]),.i2(intermediate_wire_4[30]),.o(intermediate_reg_4[15])); 
xor_module xor_module_inst_4_84(.clk(clk),.reset(reset),.i1(intermediate_wire_4[29]),.i2(intermediate_wire_4[28]),.o(intermediate_reg_4[14])); 
xor_module xor_module_inst_4_85(.clk(clk),.reset(reset),.i1(intermediate_wire_4[27]),.i2(intermediate_wire_4[26]),.o(intermediate_reg_4[13])); 
fsm fsm_inst_4_86(.clk(clk),.reset(reset),.i1(intermediate_wire_4[25]),.i2(intermediate_wire_4[24]),.o(intermediate_reg_4[12])); 
xor_module xor_module_inst_4_87(.clk(clk),.reset(reset),.i1(intermediate_wire_4[23]),.i2(intermediate_wire_4[22]),.o(intermediate_reg_4[11])); 
xor_module xor_module_inst_4_88(.clk(clk),.reset(reset),.i1(intermediate_wire_4[21]),.i2(intermediate_wire_4[20]),.o(intermediate_reg_4[10])); 
fsm fsm_inst_4_89(.clk(clk),.reset(reset),.i1(intermediate_wire_4[19]),.i2(intermediate_wire_4[18]),.o(intermediate_reg_4[9])); 
xor_module xor_module_inst_4_90(.clk(clk),.reset(reset),.i1(intermediate_wire_4[17]),.i2(intermediate_wire_4[16]),.o(intermediate_reg_4[8])); 
fsm fsm_inst_4_91(.clk(clk),.reset(reset),.i1(intermediate_wire_4[15]),.i2(intermediate_wire_4[14]),.o(intermediate_reg_4[7])); 
fsm fsm_inst_4_92(.clk(clk),.reset(reset),.i1(intermediate_wire_4[13]),.i2(intermediate_wire_4[12]),.o(intermediate_reg_4[6])); 
xor_module xor_module_inst_4_93(.clk(clk),.reset(reset),.i1(intermediate_wire_4[11]),.i2(intermediate_wire_4[10]),.o(intermediate_reg_4[5])); 
xor_module xor_module_inst_4_94(.clk(clk),.reset(reset),.i1(intermediate_wire_4[9]),.i2(intermediate_wire_4[8]),.o(intermediate_reg_4[4])); 
fsm fsm_inst_4_95(.clk(clk),.reset(reset),.i1(intermediate_wire_4[7]),.i2(intermediate_wire_4[6]),.o(intermediate_reg_4[3])); 
xor_module xor_module_inst_4_96(.clk(clk),.reset(reset),.i1(intermediate_wire_4[5]),.i2(intermediate_wire_4[4]),.o(intermediate_reg_4[2])); 
xor_module xor_module_inst_4_97(.clk(clk),.reset(reset),.i1(intermediate_wire_4[3]),.i2(intermediate_wire_4[2]),.o(intermediate_reg_4[1])); 
xor_module xor_module_inst_4_98(.clk(clk),.reset(reset),.i1(intermediate_wire_4[1]),.i2(intermediate_wire_4[0]),.o(intermediate_reg_4[0])); 
wire [97:0]intermediate_wire_5; 
assign intermediate_wire_5[97] = intermediate_reg_4[98]^intermediate_reg_4[97] ; 
assign intermediate_wire_5[96:0] = intermediate_reg_4[96:0] ; 
always@(posedge clk) begin 
outp [97:0] <= intermediate_wire_5; 
outp[171:98] <= intermediate_wire_5[73:0] ; 
end 
endmodule 
 

module interface_12(input [2207:0] inp, output reg [2367:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[2207:0] <= inp ; 
outp[2367:2208] <= inp[159:0] ; 
end 
endmodule 

module interface_14(input [250:0] inp, output reg [2015:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[250:0] <= inp ; 
outp[501:251] <= inp ; 
outp[752:502] <= inp ; 
outp[1003:753] <= inp ; 
outp[1254:1004] <= inp ; 
outp[1505:1255] <= inp ; 
outp[1756:1506] <= inp ; 
outp[2007:1757] <= inp ; 
outp[2015:2008] <= inp[7:0] ; 
end 
endmodule 

module interface_15(input [3075:0] inp, output reg [3699:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[3075:0] <= inp ; 
outp[3699:3076] <= inp[623:0] ; 
end 
endmodule 

module interface_16(input [1220:0] inp, output reg [257:0] outp, input clk, input reset);
reg [1220:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
wire [1219:0]intermediate_wire_1; 
assign intermediate_wire_1[1219] = intermediate_reg_0[1220]^intermediate_reg_0[1219] ; 
assign intermediate_wire_1[1218:0] = intermediate_reg_0[1218:0] ; 
reg [609:0]intermediate_reg_1; 
 
fsm fsm_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
xor_module xor_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
xor_module xor_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
fsm fsm_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
fsm fsm_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
fsm fsm_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
xor_module xor_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
fsm fsm_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
fsm fsm_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
xor_module xor_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
fsm fsm_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
fsm fsm_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
xor_module xor_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
fsm fsm_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
xor_module xor_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
xor_module xor_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
fsm fsm_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
fsm fsm_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
fsm fsm_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
fsm fsm_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
fsm fsm_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
fsm fsm_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
xor_module xor_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
fsm fsm_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
xor_module xor_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
fsm fsm_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
xor_module xor_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
fsm fsm_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
fsm fsm_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
fsm fsm_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
fsm fsm_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
xor_module xor_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
xor_module xor_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
xor_module xor_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
xor_module xor_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
fsm fsm_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
xor_module xor_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
fsm fsm_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
xor_module xor_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
fsm fsm_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
fsm fsm_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
xor_module xor_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
fsm fsm_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
fsm fsm_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
fsm fsm_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
fsm fsm_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
fsm fsm_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
fsm fsm_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
fsm fsm_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
fsm fsm_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
fsm fsm_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
fsm fsm_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
fsm fsm_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
fsm fsm_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
fsm fsm_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
xor_module xor_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
fsm fsm_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
xor_module xor_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
fsm fsm_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
fsm fsm_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
fsm fsm_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
xor_module xor_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
xor_module xor_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
fsm fsm_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
xor_module xor_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
fsm fsm_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
fsm fsm_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
xor_module xor_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
fsm fsm_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
fsm fsm_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
fsm fsm_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
xor_module xor_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
fsm fsm_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
xor_module xor_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
fsm fsm_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
fsm fsm_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
fsm fsm_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
xor_module xor_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
fsm fsm_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
fsm fsm_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
fsm fsm_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
fsm fsm_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
xor_module xor_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
fsm fsm_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
fsm fsm_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
fsm fsm_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
fsm fsm_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
fsm fsm_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
fsm fsm_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
fsm fsm_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
fsm fsm_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
fsm fsm_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
fsm fsm_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
xor_module xor_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
fsm fsm_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
xor_module xor_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
fsm fsm_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
fsm fsm_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
fsm fsm_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
fsm fsm_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
xor_module xor_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
fsm fsm_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
xor_module xor_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
xor_module xor_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
fsm fsm_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
fsm fsm_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
fsm fsm_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
fsm fsm_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
xor_module xor_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
fsm fsm_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
xor_module xor_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
fsm fsm_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
xor_module xor_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
fsm fsm_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
fsm fsm_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
fsm fsm_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
xor_module xor_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
xor_module xor_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
fsm fsm_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
fsm fsm_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
xor_module xor_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
fsm fsm_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
fsm fsm_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
fsm fsm_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
xor_module xor_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
fsm fsm_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
xor_module xor_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
xor_module xor_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
xor_module xor_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
fsm fsm_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
fsm fsm_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
fsm fsm_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
fsm fsm_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
xor_module xor_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
xor_module xor_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
fsm fsm_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
fsm fsm_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
fsm fsm_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
xor_module xor_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
fsm fsm_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
xor_module xor_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
fsm fsm_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
fsm fsm_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
fsm fsm_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
fsm fsm_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
fsm fsm_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
xor_module xor_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
fsm fsm_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
xor_module xor_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
xor_module xor_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
fsm fsm_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
fsm fsm_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
fsm fsm_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
fsm fsm_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
fsm fsm_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
fsm fsm_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
fsm fsm_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
fsm fsm_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
fsm fsm_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
fsm fsm_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
xor_module xor_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
xor_module xor_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
fsm fsm_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
fsm fsm_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
fsm fsm_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
fsm fsm_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
fsm fsm_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
xor_module xor_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
fsm fsm_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
fsm fsm_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
fsm fsm_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
fsm fsm_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
fsm fsm_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
fsm fsm_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
fsm fsm_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
fsm fsm_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
fsm fsm_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
fsm fsm_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
xor_module xor_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
fsm fsm_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
fsm fsm_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
fsm fsm_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
fsm fsm_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
fsm fsm_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
fsm fsm_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
fsm fsm_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
xor_module xor_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
fsm fsm_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
fsm fsm_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
fsm fsm_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
fsm fsm_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
xor_module xor_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
fsm fsm_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
xor_module xor_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
fsm fsm_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
xor_module xor_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
fsm fsm_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
xor_module xor_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
xor_module xor_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
fsm fsm_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
fsm fsm_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
fsm fsm_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
fsm fsm_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
fsm fsm_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
fsm fsm_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
fsm fsm_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
fsm fsm_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
fsm fsm_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
fsm fsm_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
fsm fsm_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
fsm fsm_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
fsm fsm_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
fsm fsm_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
fsm fsm_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
fsm fsm_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
fsm fsm_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
fsm fsm_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
fsm fsm_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
fsm fsm_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
xor_module xor_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
xor_module xor_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
xor_module xor_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
xor_module xor_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
fsm fsm_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
xor_module xor_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
xor_module xor_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
fsm fsm_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
fsm fsm_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
xor_module xor_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
fsm fsm_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
xor_module xor_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
xor_module xor_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
fsm fsm_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
fsm fsm_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
fsm fsm_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
fsm fsm_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
fsm fsm_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
fsm fsm_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
fsm fsm_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
fsm fsm_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
xor_module xor_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
xor_module xor_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
xor_module xor_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
fsm fsm_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
fsm fsm_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
xor_module xor_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
xor_module xor_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
fsm fsm_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
fsm fsm_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
fsm fsm_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
fsm fsm_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
xor_module xor_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
xor_module xor_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
fsm fsm_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
fsm fsm_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
fsm fsm_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
xor_module xor_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
fsm fsm_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
fsm fsm_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
fsm fsm_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
xor_module xor_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
fsm fsm_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
xor_module xor_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
xor_module xor_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
xor_module xor_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
fsm fsm_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
fsm fsm_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
fsm fsm_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
xor_module xor_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
fsm fsm_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
fsm fsm_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
xor_module xor_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
fsm fsm_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
xor_module xor_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
fsm fsm_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
fsm fsm_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
fsm fsm_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
fsm fsm_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
fsm fsm_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
fsm fsm_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
xor_module xor_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
xor_module xor_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
xor_module xor_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
xor_module xor_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
fsm fsm_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
fsm fsm_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
fsm fsm_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
xor_module xor_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
xor_module xor_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
xor_module xor_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
xor_module xor_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
xor_module xor_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
fsm fsm_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
xor_module xor_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
fsm fsm_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
fsm fsm_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
fsm fsm_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
xor_module xor_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
fsm fsm_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
fsm fsm_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
xor_module xor_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
fsm fsm_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
fsm fsm_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
fsm fsm_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
fsm fsm_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
fsm fsm_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
fsm fsm_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
fsm fsm_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
xor_module xor_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
xor_module xor_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
fsm fsm_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
fsm fsm_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
fsm fsm_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
fsm fsm_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
fsm fsm_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
fsm fsm_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
fsm fsm_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
fsm fsm_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
fsm fsm_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
fsm fsm_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
xor_module xor_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
fsm fsm_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
xor_module xor_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
xor_module xor_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
xor_module xor_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
xor_module xor_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
fsm fsm_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
fsm fsm_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
fsm fsm_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
xor_module xor_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
fsm fsm_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
fsm fsm_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
fsm fsm_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
fsm fsm_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
fsm fsm_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
xor_module xor_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
xor_module xor_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
xor_module xor_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
fsm fsm_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
xor_module xor_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
fsm fsm_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
reg [304:0]intermediate_reg_2; 
 
fsm fsm_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304])); 
fsm fsm_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
fsm fsm_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302])); 
fsm fsm_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
xor_module xor_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300])); 
xor_module xor_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299])); 
fsm fsm_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298])); 
xor_module xor_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297])); 
xor_module xor_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
fsm fsm_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
fsm fsm_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294])); 
fsm fsm_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
xor_module xor_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292])); 
fsm fsm_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291])); 
xor_module xor_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290])); 
xor_module xor_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289])); 
xor_module xor_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288])); 
xor_module xor_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287])); 
xor_module xor_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286])); 
fsm fsm_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
xor_module xor_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284])); 
fsm fsm_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
xor_module xor_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282])); 
xor_module xor_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281])); 
fsm fsm_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280])); 
xor_module xor_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279])); 
fsm fsm_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278])); 
xor_module xor_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277])); 
xor_module xor_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276])); 
xor_module xor_module_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275])); 
fsm fsm_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
fsm fsm_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
xor_module xor_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
xor_module xor_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
fsm fsm_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270])); 
xor_module xor_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
fsm fsm_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268])); 
fsm fsm_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267])); 
xor_module xor_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266])); 
xor_module xor_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
fsm fsm_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264])); 
xor_module xor_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263])); 
fsm fsm_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
xor_module xor_module_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261])); 
xor_module xor_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
fsm fsm_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259])); 
xor_module xor_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258])); 
xor_module xor_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257])); 
xor_module xor_module_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
fsm fsm_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255])); 
fsm fsm_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254])); 
fsm fsm_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253])); 
fsm fsm_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252])); 
fsm fsm_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
fsm fsm_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250])); 
xor_module xor_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
fsm fsm_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248])); 
xor_module xor_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247])); 
xor_module xor_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246])); 
fsm fsm_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
xor_module xor_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244])); 
xor_module xor_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243])); 
fsm fsm_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242])); 
fsm fsm_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
fsm fsm_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240])); 
xor_module xor_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239])); 
xor_module xor_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
xor_module xor_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
fsm fsm_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236])); 
fsm fsm_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235])); 
xor_module xor_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
fsm fsm_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233])); 
xor_module xor_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232])); 
fsm fsm_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231])); 
fsm fsm_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230])); 
fsm fsm_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229])); 
fsm fsm_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
fsm fsm_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227])); 
xor_module xor_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
xor_module xor_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
xor_module xor_module_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224])); 
fsm fsm_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223])); 
fsm fsm_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
fsm fsm_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221])); 
fsm fsm_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220])); 
xor_module xor_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219])); 
fsm fsm_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
fsm fsm_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217])); 
xor_module xor_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216])); 
fsm fsm_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215])); 
xor_module xor_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214])); 
fsm fsm_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
xor_module xor_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
fsm fsm_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
xor_module xor_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
fsm fsm_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209])); 
xor_module xor_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208])); 
xor_module xor_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
xor_module xor_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
fsm fsm_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
fsm fsm_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204])); 
xor_module xor_module_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203])); 
xor_module xor_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202])); 
xor_module xor_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201])); 
fsm fsm_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200])); 
xor_module xor_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
xor_module xor_module_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198])); 
xor_module xor_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197])); 
xor_module xor_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
xor_module xor_module_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195])); 
xor_module xor_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194])); 
xor_module xor_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193])); 
xor_module xor_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
xor_module xor_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
fsm fsm_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190])); 
fsm fsm_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189])); 
fsm fsm_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
fsm fsm_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
fsm fsm_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186])); 
xor_module xor_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185])); 
fsm fsm_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
fsm fsm_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183])); 
fsm fsm_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182])); 
fsm fsm_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181])); 
fsm fsm_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180])); 
fsm fsm_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179])); 
fsm fsm_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178])); 
fsm fsm_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
xor_module xor_module_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176])); 
fsm fsm_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175])); 
xor_module xor_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174])); 
xor_module xor_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
fsm fsm_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
xor_module xor_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
fsm fsm_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
fsm fsm_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169])); 
xor_module xor_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168])); 
fsm fsm_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167])); 
fsm fsm_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166])); 
fsm fsm_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
fsm fsm_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164])); 
xor_module xor_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
xor_module xor_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162])); 
xor_module xor_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161])); 
fsm fsm_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160])); 
fsm fsm_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
fsm fsm_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158])); 
fsm fsm_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157])); 
xor_module xor_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156])); 
xor_module xor_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155])); 
fsm fsm_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154])); 
fsm fsm_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153])); 
fsm fsm_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152])); 
fsm fsm_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151])); 
fsm fsm_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
fsm fsm_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
fsm fsm_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148])); 
fsm fsm_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147])); 
fsm fsm_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146])); 
xor_module xor_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145])); 
fsm fsm_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144])); 
xor_module xor_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143])); 
fsm fsm_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142])); 
fsm fsm_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141])); 
xor_module xor_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140])); 
fsm fsm_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139])); 
fsm fsm_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138])); 
xor_module xor_module_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
xor_module xor_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136])); 
xor_module xor_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135])); 
xor_module xor_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
xor_module xor_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133])); 
xor_module xor_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132])); 
xor_module xor_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131])); 
fsm fsm_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130])); 
xor_module xor_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129])); 
xor_module xor_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
fsm fsm_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
xor_module xor_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126])); 
fsm fsm_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
fsm fsm_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124])); 
fsm fsm_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123])); 
fsm fsm_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
fsm fsm_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121])); 
fsm fsm_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120])); 
xor_module xor_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119])); 
xor_module xor_module_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118])); 
xor_module xor_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117])); 
fsm fsm_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116])); 
fsm fsm_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115])); 
xor_module xor_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
fsm fsm_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113])); 
xor_module xor_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
fsm fsm_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111])); 
fsm fsm_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
xor_module xor_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
xor_module xor_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
fsm fsm_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107])); 
xor_module xor_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
xor_module xor_module_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105])); 
fsm fsm_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104])); 
fsm fsm_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
fsm fsm_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102])); 
xor_module xor_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
xor_module xor_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100])); 
fsm fsm_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99])); 
xor_module xor_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98])); 
xor_module xor_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
fsm fsm_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96])); 
xor_module xor_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95])); 
fsm fsm_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94])); 
fsm fsm_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
fsm fsm_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92])); 
fsm fsm_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91])); 
xor_module xor_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
xor_module xor_module_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89])); 
fsm fsm_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88])); 
xor_module xor_module_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
fsm fsm_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
fsm fsm_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
xor_module xor_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
xor_module xor_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
fsm fsm_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82])); 
fsm fsm_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
xor_module xor_module_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80])); 
xor_module xor_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79])); 
fsm fsm_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78])); 
fsm fsm_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
fsm fsm_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76])); 
fsm fsm_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
xor_module xor_module_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74])); 
xor_module xor_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73])); 
xor_module xor_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72])); 
xor_module xor_module_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71])); 
xor_module xor_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
xor_module xor_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69])); 
xor_module xor_module_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68])); 
fsm fsm_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67])); 
xor_module xor_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66])); 
xor_module xor_module_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65])); 
fsm fsm_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64])); 
xor_module xor_module_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
xor_module xor_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
xor_module xor_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
xor_module xor_module_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60])); 
xor_module xor_module_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59])); 
xor_module xor_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
xor_module xor_module_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57])); 
xor_module xor_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56])); 
xor_module xor_module_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55])); 
xor_module xor_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54])); 
fsm fsm_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
fsm fsm_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
xor_module xor_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51])); 
fsm fsm_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
fsm fsm_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
xor_module xor_module_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48])); 
fsm fsm_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47])); 
xor_module xor_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46])); 
fsm fsm_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45])); 
xor_module xor_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44])); 
xor_module xor_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
xor_module xor_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42])); 
fsm fsm_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
fsm fsm_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40])); 
fsm fsm_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39])); 
xor_module xor_module_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38])); 
xor_module xor_module_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
xor_module xor_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36])); 
xor_module xor_module_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35])); 
xor_module xor_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34])); 
xor_module xor_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33])); 
xor_module xor_module_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32])); 
xor_module xor_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
xor_module xor_module_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
xor_module xor_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29])); 
fsm fsm_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
xor_module xor_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27])); 
fsm fsm_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26])); 
xor_module xor_module_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25])); 
fsm fsm_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
xor_module xor_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23])); 
fsm fsm_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22])); 
xor_module xor_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21])); 
fsm fsm_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20])); 
xor_module xor_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
xor_module xor_module_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18])); 
xor_module xor_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17])); 
fsm fsm_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
fsm fsm_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15])); 
xor_module xor_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14])); 
fsm fsm_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13])); 
fsm fsm_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12])); 
xor_module xor_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11])); 
xor_module xor_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10])); 
fsm fsm_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
fsm fsm_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8])); 
xor_module xor_module_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
xor_module xor_module_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6])); 
xor_module xor_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5])); 
fsm fsm_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
fsm fsm_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
xor_module xor_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2])); 
xor_module xor_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
fsm fsm_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0])); 
wire [303:0]intermediate_wire_3; 
assign intermediate_wire_3[303] = intermediate_reg_2[304]^intermediate_reg_2[303] ; 
assign intermediate_wire_3[302:0] = intermediate_reg_2[302:0] ; 
reg [151:0]intermediate_reg_3; 
 
xor_module xor_module_inst_3_0(.clk(clk),.reset(reset),.i1(intermediate_wire_3[303]),.i2(intermediate_wire_3[302]),.o(intermediate_reg_3[151])); 
xor_module xor_module_inst_3_1(.clk(clk),.reset(reset),.i1(intermediate_wire_3[301]),.i2(intermediate_wire_3[300]),.o(intermediate_reg_3[150])); 
fsm fsm_inst_3_2(.clk(clk),.reset(reset),.i1(intermediate_wire_3[299]),.i2(intermediate_wire_3[298]),.o(intermediate_reg_3[149])); 
fsm fsm_inst_3_3(.clk(clk),.reset(reset),.i1(intermediate_wire_3[297]),.i2(intermediate_wire_3[296]),.o(intermediate_reg_3[148])); 
xor_module xor_module_inst_3_4(.clk(clk),.reset(reset),.i1(intermediate_wire_3[295]),.i2(intermediate_wire_3[294]),.o(intermediate_reg_3[147])); 
fsm fsm_inst_3_5(.clk(clk),.reset(reset),.i1(intermediate_wire_3[293]),.i2(intermediate_wire_3[292]),.o(intermediate_reg_3[146])); 
xor_module xor_module_inst_3_6(.clk(clk),.reset(reset),.i1(intermediate_wire_3[291]),.i2(intermediate_wire_3[290]),.o(intermediate_reg_3[145])); 
fsm fsm_inst_3_7(.clk(clk),.reset(reset),.i1(intermediate_wire_3[289]),.i2(intermediate_wire_3[288]),.o(intermediate_reg_3[144])); 
xor_module xor_module_inst_3_8(.clk(clk),.reset(reset),.i1(intermediate_wire_3[287]),.i2(intermediate_wire_3[286]),.o(intermediate_reg_3[143])); 
fsm fsm_inst_3_9(.clk(clk),.reset(reset),.i1(intermediate_wire_3[285]),.i2(intermediate_wire_3[284]),.o(intermediate_reg_3[142])); 
xor_module xor_module_inst_3_10(.clk(clk),.reset(reset),.i1(intermediate_wire_3[283]),.i2(intermediate_wire_3[282]),.o(intermediate_reg_3[141])); 
xor_module xor_module_inst_3_11(.clk(clk),.reset(reset),.i1(intermediate_wire_3[281]),.i2(intermediate_wire_3[280]),.o(intermediate_reg_3[140])); 
xor_module xor_module_inst_3_12(.clk(clk),.reset(reset),.i1(intermediate_wire_3[279]),.i2(intermediate_wire_3[278]),.o(intermediate_reg_3[139])); 
xor_module xor_module_inst_3_13(.clk(clk),.reset(reset),.i1(intermediate_wire_3[277]),.i2(intermediate_wire_3[276]),.o(intermediate_reg_3[138])); 
fsm fsm_inst_3_14(.clk(clk),.reset(reset),.i1(intermediate_wire_3[275]),.i2(intermediate_wire_3[274]),.o(intermediate_reg_3[137])); 
xor_module xor_module_inst_3_15(.clk(clk),.reset(reset),.i1(intermediate_wire_3[273]),.i2(intermediate_wire_3[272]),.o(intermediate_reg_3[136])); 
xor_module xor_module_inst_3_16(.clk(clk),.reset(reset),.i1(intermediate_wire_3[271]),.i2(intermediate_wire_3[270]),.o(intermediate_reg_3[135])); 
xor_module xor_module_inst_3_17(.clk(clk),.reset(reset),.i1(intermediate_wire_3[269]),.i2(intermediate_wire_3[268]),.o(intermediate_reg_3[134])); 
xor_module xor_module_inst_3_18(.clk(clk),.reset(reset),.i1(intermediate_wire_3[267]),.i2(intermediate_wire_3[266]),.o(intermediate_reg_3[133])); 
xor_module xor_module_inst_3_19(.clk(clk),.reset(reset),.i1(intermediate_wire_3[265]),.i2(intermediate_wire_3[264]),.o(intermediate_reg_3[132])); 
fsm fsm_inst_3_20(.clk(clk),.reset(reset),.i1(intermediate_wire_3[263]),.i2(intermediate_wire_3[262]),.o(intermediate_reg_3[131])); 
fsm fsm_inst_3_21(.clk(clk),.reset(reset),.i1(intermediate_wire_3[261]),.i2(intermediate_wire_3[260]),.o(intermediate_reg_3[130])); 
fsm fsm_inst_3_22(.clk(clk),.reset(reset),.i1(intermediate_wire_3[259]),.i2(intermediate_wire_3[258]),.o(intermediate_reg_3[129])); 
xor_module xor_module_inst_3_23(.clk(clk),.reset(reset),.i1(intermediate_wire_3[257]),.i2(intermediate_wire_3[256]),.o(intermediate_reg_3[128])); 
fsm fsm_inst_3_24(.clk(clk),.reset(reset),.i1(intermediate_wire_3[255]),.i2(intermediate_wire_3[254]),.o(intermediate_reg_3[127])); 
xor_module xor_module_inst_3_25(.clk(clk),.reset(reset),.i1(intermediate_wire_3[253]),.i2(intermediate_wire_3[252]),.o(intermediate_reg_3[126])); 
xor_module xor_module_inst_3_26(.clk(clk),.reset(reset),.i1(intermediate_wire_3[251]),.i2(intermediate_wire_3[250]),.o(intermediate_reg_3[125])); 
xor_module xor_module_inst_3_27(.clk(clk),.reset(reset),.i1(intermediate_wire_3[249]),.i2(intermediate_wire_3[248]),.o(intermediate_reg_3[124])); 
xor_module xor_module_inst_3_28(.clk(clk),.reset(reset),.i1(intermediate_wire_3[247]),.i2(intermediate_wire_3[246]),.o(intermediate_reg_3[123])); 
xor_module xor_module_inst_3_29(.clk(clk),.reset(reset),.i1(intermediate_wire_3[245]),.i2(intermediate_wire_3[244]),.o(intermediate_reg_3[122])); 
xor_module xor_module_inst_3_30(.clk(clk),.reset(reset),.i1(intermediate_wire_3[243]),.i2(intermediate_wire_3[242]),.o(intermediate_reg_3[121])); 
fsm fsm_inst_3_31(.clk(clk),.reset(reset),.i1(intermediate_wire_3[241]),.i2(intermediate_wire_3[240]),.o(intermediate_reg_3[120])); 
xor_module xor_module_inst_3_32(.clk(clk),.reset(reset),.i1(intermediate_wire_3[239]),.i2(intermediate_wire_3[238]),.o(intermediate_reg_3[119])); 
xor_module xor_module_inst_3_33(.clk(clk),.reset(reset),.i1(intermediate_wire_3[237]),.i2(intermediate_wire_3[236]),.o(intermediate_reg_3[118])); 
xor_module xor_module_inst_3_34(.clk(clk),.reset(reset),.i1(intermediate_wire_3[235]),.i2(intermediate_wire_3[234]),.o(intermediate_reg_3[117])); 
xor_module xor_module_inst_3_35(.clk(clk),.reset(reset),.i1(intermediate_wire_3[233]),.i2(intermediate_wire_3[232]),.o(intermediate_reg_3[116])); 
fsm fsm_inst_3_36(.clk(clk),.reset(reset),.i1(intermediate_wire_3[231]),.i2(intermediate_wire_3[230]),.o(intermediate_reg_3[115])); 
xor_module xor_module_inst_3_37(.clk(clk),.reset(reset),.i1(intermediate_wire_3[229]),.i2(intermediate_wire_3[228]),.o(intermediate_reg_3[114])); 
xor_module xor_module_inst_3_38(.clk(clk),.reset(reset),.i1(intermediate_wire_3[227]),.i2(intermediate_wire_3[226]),.o(intermediate_reg_3[113])); 
fsm fsm_inst_3_39(.clk(clk),.reset(reset),.i1(intermediate_wire_3[225]),.i2(intermediate_wire_3[224]),.o(intermediate_reg_3[112])); 
fsm fsm_inst_3_40(.clk(clk),.reset(reset),.i1(intermediate_wire_3[223]),.i2(intermediate_wire_3[222]),.o(intermediate_reg_3[111])); 
fsm fsm_inst_3_41(.clk(clk),.reset(reset),.i1(intermediate_wire_3[221]),.i2(intermediate_wire_3[220]),.o(intermediate_reg_3[110])); 
fsm fsm_inst_3_42(.clk(clk),.reset(reset),.i1(intermediate_wire_3[219]),.i2(intermediate_wire_3[218]),.o(intermediate_reg_3[109])); 
fsm fsm_inst_3_43(.clk(clk),.reset(reset),.i1(intermediate_wire_3[217]),.i2(intermediate_wire_3[216]),.o(intermediate_reg_3[108])); 
xor_module xor_module_inst_3_44(.clk(clk),.reset(reset),.i1(intermediate_wire_3[215]),.i2(intermediate_wire_3[214]),.o(intermediate_reg_3[107])); 
xor_module xor_module_inst_3_45(.clk(clk),.reset(reset),.i1(intermediate_wire_3[213]),.i2(intermediate_wire_3[212]),.o(intermediate_reg_3[106])); 
xor_module xor_module_inst_3_46(.clk(clk),.reset(reset),.i1(intermediate_wire_3[211]),.i2(intermediate_wire_3[210]),.o(intermediate_reg_3[105])); 
xor_module xor_module_inst_3_47(.clk(clk),.reset(reset),.i1(intermediate_wire_3[209]),.i2(intermediate_wire_3[208]),.o(intermediate_reg_3[104])); 
fsm fsm_inst_3_48(.clk(clk),.reset(reset),.i1(intermediate_wire_3[207]),.i2(intermediate_wire_3[206]),.o(intermediate_reg_3[103])); 
xor_module xor_module_inst_3_49(.clk(clk),.reset(reset),.i1(intermediate_wire_3[205]),.i2(intermediate_wire_3[204]),.o(intermediate_reg_3[102])); 
xor_module xor_module_inst_3_50(.clk(clk),.reset(reset),.i1(intermediate_wire_3[203]),.i2(intermediate_wire_3[202]),.o(intermediate_reg_3[101])); 
xor_module xor_module_inst_3_51(.clk(clk),.reset(reset),.i1(intermediate_wire_3[201]),.i2(intermediate_wire_3[200]),.o(intermediate_reg_3[100])); 
xor_module xor_module_inst_3_52(.clk(clk),.reset(reset),.i1(intermediate_wire_3[199]),.i2(intermediate_wire_3[198]),.o(intermediate_reg_3[99])); 
xor_module xor_module_inst_3_53(.clk(clk),.reset(reset),.i1(intermediate_wire_3[197]),.i2(intermediate_wire_3[196]),.o(intermediate_reg_3[98])); 
fsm fsm_inst_3_54(.clk(clk),.reset(reset),.i1(intermediate_wire_3[195]),.i2(intermediate_wire_3[194]),.o(intermediate_reg_3[97])); 
xor_module xor_module_inst_3_55(.clk(clk),.reset(reset),.i1(intermediate_wire_3[193]),.i2(intermediate_wire_3[192]),.o(intermediate_reg_3[96])); 
fsm fsm_inst_3_56(.clk(clk),.reset(reset),.i1(intermediate_wire_3[191]),.i2(intermediate_wire_3[190]),.o(intermediate_reg_3[95])); 
fsm fsm_inst_3_57(.clk(clk),.reset(reset),.i1(intermediate_wire_3[189]),.i2(intermediate_wire_3[188]),.o(intermediate_reg_3[94])); 
xor_module xor_module_inst_3_58(.clk(clk),.reset(reset),.i1(intermediate_wire_3[187]),.i2(intermediate_wire_3[186]),.o(intermediate_reg_3[93])); 
fsm fsm_inst_3_59(.clk(clk),.reset(reset),.i1(intermediate_wire_3[185]),.i2(intermediate_wire_3[184]),.o(intermediate_reg_3[92])); 
fsm fsm_inst_3_60(.clk(clk),.reset(reset),.i1(intermediate_wire_3[183]),.i2(intermediate_wire_3[182]),.o(intermediate_reg_3[91])); 
fsm fsm_inst_3_61(.clk(clk),.reset(reset),.i1(intermediate_wire_3[181]),.i2(intermediate_wire_3[180]),.o(intermediate_reg_3[90])); 
xor_module xor_module_inst_3_62(.clk(clk),.reset(reset),.i1(intermediate_wire_3[179]),.i2(intermediate_wire_3[178]),.o(intermediate_reg_3[89])); 
fsm fsm_inst_3_63(.clk(clk),.reset(reset),.i1(intermediate_wire_3[177]),.i2(intermediate_wire_3[176]),.o(intermediate_reg_3[88])); 
xor_module xor_module_inst_3_64(.clk(clk),.reset(reset),.i1(intermediate_wire_3[175]),.i2(intermediate_wire_3[174]),.o(intermediate_reg_3[87])); 
fsm fsm_inst_3_65(.clk(clk),.reset(reset),.i1(intermediate_wire_3[173]),.i2(intermediate_wire_3[172]),.o(intermediate_reg_3[86])); 
fsm fsm_inst_3_66(.clk(clk),.reset(reset),.i1(intermediate_wire_3[171]),.i2(intermediate_wire_3[170]),.o(intermediate_reg_3[85])); 
xor_module xor_module_inst_3_67(.clk(clk),.reset(reset),.i1(intermediate_wire_3[169]),.i2(intermediate_wire_3[168]),.o(intermediate_reg_3[84])); 
fsm fsm_inst_3_68(.clk(clk),.reset(reset),.i1(intermediate_wire_3[167]),.i2(intermediate_wire_3[166]),.o(intermediate_reg_3[83])); 
fsm fsm_inst_3_69(.clk(clk),.reset(reset),.i1(intermediate_wire_3[165]),.i2(intermediate_wire_3[164]),.o(intermediate_reg_3[82])); 
fsm fsm_inst_3_70(.clk(clk),.reset(reset),.i1(intermediate_wire_3[163]),.i2(intermediate_wire_3[162]),.o(intermediate_reg_3[81])); 
fsm fsm_inst_3_71(.clk(clk),.reset(reset),.i1(intermediate_wire_3[161]),.i2(intermediate_wire_3[160]),.o(intermediate_reg_3[80])); 
fsm fsm_inst_3_72(.clk(clk),.reset(reset),.i1(intermediate_wire_3[159]),.i2(intermediate_wire_3[158]),.o(intermediate_reg_3[79])); 
xor_module xor_module_inst_3_73(.clk(clk),.reset(reset),.i1(intermediate_wire_3[157]),.i2(intermediate_wire_3[156]),.o(intermediate_reg_3[78])); 
xor_module xor_module_inst_3_74(.clk(clk),.reset(reset),.i1(intermediate_wire_3[155]),.i2(intermediate_wire_3[154]),.o(intermediate_reg_3[77])); 
xor_module xor_module_inst_3_75(.clk(clk),.reset(reset),.i1(intermediate_wire_3[153]),.i2(intermediate_wire_3[152]),.o(intermediate_reg_3[76])); 
fsm fsm_inst_3_76(.clk(clk),.reset(reset),.i1(intermediate_wire_3[151]),.i2(intermediate_wire_3[150]),.o(intermediate_reg_3[75])); 
xor_module xor_module_inst_3_77(.clk(clk),.reset(reset),.i1(intermediate_wire_3[149]),.i2(intermediate_wire_3[148]),.o(intermediate_reg_3[74])); 
xor_module xor_module_inst_3_78(.clk(clk),.reset(reset),.i1(intermediate_wire_3[147]),.i2(intermediate_wire_3[146]),.o(intermediate_reg_3[73])); 
xor_module xor_module_inst_3_79(.clk(clk),.reset(reset),.i1(intermediate_wire_3[145]),.i2(intermediate_wire_3[144]),.o(intermediate_reg_3[72])); 
fsm fsm_inst_3_80(.clk(clk),.reset(reset),.i1(intermediate_wire_3[143]),.i2(intermediate_wire_3[142]),.o(intermediate_reg_3[71])); 
fsm fsm_inst_3_81(.clk(clk),.reset(reset),.i1(intermediate_wire_3[141]),.i2(intermediate_wire_3[140]),.o(intermediate_reg_3[70])); 
xor_module xor_module_inst_3_82(.clk(clk),.reset(reset),.i1(intermediate_wire_3[139]),.i2(intermediate_wire_3[138]),.o(intermediate_reg_3[69])); 
fsm fsm_inst_3_83(.clk(clk),.reset(reset),.i1(intermediate_wire_3[137]),.i2(intermediate_wire_3[136]),.o(intermediate_reg_3[68])); 
xor_module xor_module_inst_3_84(.clk(clk),.reset(reset),.i1(intermediate_wire_3[135]),.i2(intermediate_wire_3[134]),.o(intermediate_reg_3[67])); 
fsm fsm_inst_3_85(.clk(clk),.reset(reset),.i1(intermediate_wire_3[133]),.i2(intermediate_wire_3[132]),.o(intermediate_reg_3[66])); 
fsm fsm_inst_3_86(.clk(clk),.reset(reset),.i1(intermediate_wire_3[131]),.i2(intermediate_wire_3[130]),.o(intermediate_reg_3[65])); 
xor_module xor_module_inst_3_87(.clk(clk),.reset(reset),.i1(intermediate_wire_3[129]),.i2(intermediate_wire_3[128]),.o(intermediate_reg_3[64])); 
xor_module xor_module_inst_3_88(.clk(clk),.reset(reset),.i1(intermediate_wire_3[127]),.i2(intermediate_wire_3[126]),.o(intermediate_reg_3[63])); 
fsm fsm_inst_3_89(.clk(clk),.reset(reset),.i1(intermediate_wire_3[125]),.i2(intermediate_wire_3[124]),.o(intermediate_reg_3[62])); 
xor_module xor_module_inst_3_90(.clk(clk),.reset(reset),.i1(intermediate_wire_3[123]),.i2(intermediate_wire_3[122]),.o(intermediate_reg_3[61])); 
fsm fsm_inst_3_91(.clk(clk),.reset(reset),.i1(intermediate_wire_3[121]),.i2(intermediate_wire_3[120]),.o(intermediate_reg_3[60])); 
xor_module xor_module_inst_3_92(.clk(clk),.reset(reset),.i1(intermediate_wire_3[119]),.i2(intermediate_wire_3[118]),.o(intermediate_reg_3[59])); 
xor_module xor_module_inst_3_93(.clk(clk),.reset(reset),.i1(intermediate_wire_3[117]),.i2(intermediate_wire_3[116]),.o(intermediate_reg_3[58])); 
fsm fsm_inst_3_94(.clk(clk),.reset(reset),.i1(intermediate_wire_3[115]),.i2(intermediate_wire_3[114]),.o(intermediate_reg_3[57])); 
xor_module xor_module_inst_3_95(.clk(clk),.reset(reset),.i1(intermediate_wire_3[113]),.i2(intermediate_wire_3[112]),.o(intermediate_reg_3[56])); 
fsm fsm_inst_3_96(.clk(clk),.reset(reset),.i1(intermediate_wire_3[111]),.i2(intermediate_wire_3[110]),.o(intermediate_reg_3[55])); 
fsm fsm_inst_3_97(.clk(clk),.reset(reset),.i1(intermediate_wire_3[109]),.i2(intermediate_wire_3[108]),.o(intermediate_reg_3[54])); 
fsm fsm_inst_3_98(.clk(clk),.reset(reset),.i1(intermediate_wire_3[107]),.i2(intermediate_wire_3[106]),.o(intermediate_reg_3[53])); 
fsm fsm_inst_3_99(.clk(clk),.reset(reset),.i1(intermediate_wire_3[105]),.i2(intermediate_wire_3[104]),.o(intermediate_reg_3[52])); 
fsm fsm_inst_3_100(.clk(clk),.reset(reset),.i1(intermediate_wire_3[103]),.i2(intermediate_wire_3[102]),.o(intermediate_reg_3[51])); 
xor_module xor_module_inst_3_101(.clk(clk),.reset(reset),.i1(intermediate_wire_3[101]),.i2(intermediate_wire_3[100]),.o(intermediate_reg_3[50])); 
xor_module xor_module_inst_3_102(.clk(clk),.reset(reset),.i1(intermediate_wire_3[99]),.i2(intermediate_wire_3[98]),.o(intermediate_reg_3[49])); 
fsm fsm_inst_3_103(.clk(clk),.reset(reset),.i1(intermediate_wire_3[97]),.i2(intermediate_wire_3[96]),.o(intermediate_reg_3[48])); 
fsm fsm_inst_3_104(.clk(clk),.reset(reset),.i1(intermediate_wire_3[95]),.i2(intermediate_wire_3[94]),.o(intermediate_reg_3[47])); 
fsm fsm_inst_3_105(.clk(clk),.reset(reset),.i1(intermediate_wire_3[93]),.i2(intermediate_wire_3[92]),.o(intermediate_reg_3[46])); 
xor_module xor_module_inst_3_106(.clk(clk),.reset(reset),.i1(intermediate_wire_3[91]),.i2(intermediate_wire_3[90]),.o(intermediate_reg_3[45])); 
fsm fsm_inst_3_107(.clk(clk),.reset(reset),.i1(intermediate_wire_3[89]),.i2(intermediate_wire_3[88]),.o(intermediate_reg_3[44])); 
fsm fsm_inst_3_108(.clk(clk),.reset(reset),.i1(intermediate_wire_3[87]),.i2(intermediate_wire_3[86]),.o(intermediate_reg_3[43])); 
xor_module xor_module_inst_3_109(.clk(clk),.reset(reset),.i1(intermediate_wire_3[85]),.i2(intermediate_wire_3[84]),.o(intermediate_reg_3[42])); 
fsm fsm_inst_3_110(.clk(clk),.reset(reset),.i1(intermediate_wire_3[83]),.i2(intermediate_wire_3[82]),.o(intermediate_reg_3[41])); 
fsm fsm_inst_3_111(.clk(clk),.reset(reset),.i1(intermediate_wire_3[81]),.i2(intermediate_wire_3[80]),.o(intermediate_reg_3[40])); 
fsm fsm_inst_3_112(.clk(clk),.reset(reset),.i1(intermediate_wire_3[79]),.i2(intermediate_wire_3[78]),.o(intermediate_reg_3[39])); 
fsm fsm_inst_3_113(.clk(clk),.reset(reset),.i1(intermediate_wire_3[77]),.i2(intermediate_wire_3[76]),.o(intermediate_reg_3[38])); 
fsm fsm_inst_3_114(.clk(clk),.reset(reset),.i1(intermediate_wire_3[75]),.i2(intermediate_wire_3[74]),.o(intermediate_reg_3[37])); 
xor_module xor_module_inst_3_115(.clk(clk),.reset(reset),.i1(intermediate_wire_3[73]),.i2(intermediate_wire_3[72]),.o(intermediate_reg_3[36])); 
fsm fsm_inst_3_116(.clk(clk),.reset(reset),.i1(intermediate_wire_3[71]),.i2(intermediate_wire_3[70]),.o(intermediate_reg_3[35])); 
xor_module xor_module_inst_3_117(.clk(clk),.reset(reset),.i1(intermediate_wire_3[69]),.i2(intermediate_wire_3[68]),.o(intermediate_reg_3[34])); 
xor_module xor_module_inst_3_118(.clk(clk),.reset(reset),.i1(intermediate_wire_3[67]),.i2(intermediate_wire_3[66]),.o(intermediate_reg_3[33])); 
fsm fsm_inst_3_119(.clk(clk),.reset(reset),.i1(intermediate_wire_3[65]),.i2(intermediate_wire_3[64]),.o(intermediate_reg_3[32])); 
xor_module xor_module_inst_3_120(.clk(clk),.reset(reset),.i1(intermediate_wire_3[63]),.i2(intermediate_wire_3[62]),.o(intermediate_reg_3[31])); 
xor_module xor_module_inst_3_121(.clk(clk),.reset(reset),.i1(intermediate_wire_3[61]),.i2(intermediate_wire_3[60]),.o(intermediate_reg_3[30])); 
fsm fsm_inst_3_122(.clk(clk),.reset(reset),.i1(intermediate_wire_3[59]),.i2(intermediate_wire_3[58]),.o(intermediate_reg_3[29])); 
fsm fsm_inst_3_123(.clk(clk),.reset(reset),.i1(intermediate_wire_3[57]),.i2(intermediate_wire_3[56]),.o(intermediate_reg_3[28])); 
fsm fsm_inst_3_124(.clk(clk),.reset(reset),.i1(intermediate_wire_3[55]),.i2(intermediate_wire_3[54]),.o(intermediate_reg_3[27])); 
xor_module xor_module_inst_3_125(.clk(clk),.reset(reset),.i1(intermediate_wire_3[53]),.i2(intermediate_wire_3[52]),.o(intermediate_reg_3[26])); 
xor_module xor_module_inst_3_126(.clk(clk),.reset(reset),.i1(intermediate_wire_3[51]),.i2(intermediate_wire_3[50]),.o(intermediate_reg_3[25])); 
fsm fsm_inst_3_127(.clk(clk),.reset(reset),.i1(intermediate_wire_3[49]),.i2(intermediate_wire_3[48]),.o(intermediate_reg_3[24])); 
fsm fsm_inst_3_128(.clk(clk),.reset(reset),.i1(intermediate_wire_3[47]),.i2(intermediate_wire_3[46]),.o(intermediate_reg_3[23])); 
xor_module xor_module_inst_3_129(.clk(clk),.reset(reset),.i1(intermediate_wire_3[45]),.i2(intermediate_wire_3[44]),.o(intermediate_reg_3[22])); 
fsm fsm_inst_3_130(.clk(clk),.reset(reset),.i1(intermediate_wire_3[43]),.i2(intermediate_wire_3[42]),.o(intermediate_reg_3[21])); 
xor_module xor_module_inst_3_131(.clk(clk),.reset(reset),.i1(intermediate_wire_3[41]),.i2(intermediate_wire_3[40]),.o(intermediate_reg_3[20])); 
xor_module xor_module_inst_3_132(.clk(clk),.reset(reset),.i1(intermediate_wire_3[39]),.i2(intermediate_wire_3[38]),.o(intermediate_reg_3[19])); 
xor_module xor_module_inst_3_133(.clk(clk),.reset(reset),.i1(intermediate_wire_3[37]),.i2(intermediate_wire_3[36]),.o(intermediate_reg_3[18])); 
fsm fsm_inst_3_134(.clk(clk),.reset(reset),.i1(intermediate_wire_3[35]),.i2(intermediate_wire_3[34]),.o(intermediate_reg_3[17])); 
fsm fsm_inst_3_135(.clk(clk),.reset(reset),.i1(intermediate_wire_3[33]),.i2(intermediate_wire_3[32]),.o(intermediate_reg_3[16])); 
xor_module xor_module_inst_3_136(.clk(clk),.reset(reset),.i1(intermediate_wire_3[31]),.i2(intermediate_wire_3[30]),.o(intermediate_reg_3[15])); 
xor_module xor_module_inst_3_137(.clk(clk),.reset(reset),.i1(intermediate_wire_3[29]),.i2(intermediate_wire_3[28]),.o(intermediate_reg_3[14])); 
xor_module xor_module_inst_3_138(.clk(clk),.reset(reset),.i1(intermediate_wire_3[27]),.i2(intermediate_wire_3[26]),.o(intermediate_reg_3[13])); 
fsm fsm_inst_3_139(.clk(clk),.reset(reset),.i1(intermediate_wire_3[25]),.i2(intermediate_wire_3[24]),.o(intermediate_reg_3[12])); 
fsm fsm_inst_3_140(.clk(clk),.reset(reset),.i1(intermediate_wire_3[23]),.i2(intermediate_wire_3[22]),.o(intermediate_reg_3[11])); 
fsm fsm_inst_3_141(.clk(clk),.reset(reset),.i1(intermediate_wire_3[21]),.i2(intermediate_wire_3[20]),.o(intermediate_reg_3[10])); 
xor_module xor_module_inst_3_142(.clk(clk),.reset(reset),.i1(intermediate_wire_3[19]),.i2(intermediate_wire_3[18]),.o(intermediate_reg_3[9])); 
fsm fsm_inst_3_143(.clk(clk),.reset(reset),.i1(intermediate_wire_3[17]),.i2(intermediate_wire_3[16]),.o(intermediate_reg_3[8])); 
xor_module xor_module_inst_3_144(.clk(clk),.reset(reset),.i1(intermediate_wire_3[15]),.i2(intermediate_wire_3[14]),.o(intermediate_reg_3[7])); 
xor_module xor_module_inst_3_145(.clk(clk),.reset(reset),.i1(intermediate_wire_3[13]),.i2(intermediate_wire_3[12]),.o(intermediate_reg_3[6])); 
fsm fsm_inst_3_146(.clk(clk),.reset(reset),.i1(intermediate_wire_3[11]),.i2(intermediate_wire_3[10]),.o(intermediate_reg_3[5])); 
fsm fsm_inst_3_147(.clk(clk),.reset(reset),.i1(intermediate_wire_3[9]),.i2(intermediate_wire_3[8]),.o(intermediate_reg_3[4])); 
xor_module xor_module_inst_3_148(.clk(clk),.reset(reset),.i1(intermediate_wire_3[7]),.i2(intermediate_wire_3[6]),.o(intermediate_reg_3[3])); 
xor_module xor_module_inst_3_149(.clk(clk),.reset(reset),.i1(intermediate_wire_3[5]),.i2(intermediate_wire_3[4]),.o(intermediate_reg_3[2])); 
fsm fsm_inst_3_150(.clk(clk),.reset(reset),.i1(intermediate_wire_3[3]),.i2(intermediate_wire_3[2]),.o(intermediate_reg_3[1])); 
xor_module xor_module_inst_3_151(.clk(clk),.reset(reset),.i1(intermediate_wire_3[1]),.i2(intermediate_wire_3[0]),.o(intermediate_reg_3[0])); 
always@(posedge clk) begin 
outp [151:0] <= intermediate_reg_3; 
outp[257:152] <= intermediate_reg_3[105:0] ; 
end 
endmodule 
 

module fifo_512_60bit_module_4(input clk, input reset, input[251:0] inp, output reg [247:0] outp); 

fifo_512_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[62:0]),.outp(outp[61:0])); 

fifo_512_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[125:63]),.outp(outp[123:62])); 

fifo_512_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[188:126]),.outp(outp[185:124])); 

fifo_512_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[251:189]),.outp(outp[247:186])); 

endmodule 

module fifo_256_40bit_module_2(input clk, input reset, input[85:0] inp, output reg [83:0] outp); 

fifo_256_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[42:0]),.outp(outp[41:0])); 

fifo_256_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[85:43]),.outp(outp[83:42])); 

endmodule 

module tensor_block_int8_module_4(input clk, input reset, input[1059:0] inp, output reg [1003:0] outp); 

tensor_block_int8_module inst_0 (.clk(clk),.reset(reset),.inp(inp[264:0]),.outp(outp[250:0])); 

tensor_block_int8_module inst_1 (.clk(clk),.reset(reset),.inp(inp[529:265]),.outp(outp[501:251])); 

tensor_block_int8_module inst_2 (.clk(clk),.reset(reset),.inp(inp[794:530]),.outp(outp[752:502])); 

tensor_block_int8_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1059:795]),.outp(outp[1003:753])); 

endmodule 

module tensor_block_int8_module_8(input clk, input reset, input[2119:0] inp, output reg [2007:0] outp); 

tensor_block_int8_module inst_0 (.clk(clk),.reset(reset),.inp(inp[264:0]),.outp(outp[250:0])); 

tensor_block_int8_module inst_1 (.clk(clk),.reset(reset),.inp(inp[529:265]),.outp(outp[501:251])); 

tensor_block_int8_module inst_2 (.clk(clk),.reset(reset),.inp(inp[794:530]),.outp(outp[752:502])); 

tensor_block_int8_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1059:795]),.outp(outp[1003:753])); 

tensor_block_int8_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1324:1060]),.outp(outp[1254:1004])); 

tensor_block_int8_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1589:1325]),.outp(outp[1505:1255])); 

tensor_block_int8_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1854:1590]),.outp(outp[1756:1506])); 

tensor_block_int8_module inst_7 (.clk(clk),.reset(reset),.inp(inp[2119:1855]),.outp(outp[2007:1757])); 

endmodule 

module dsp_chain_4_int_sop_2_module_6(input clk, input reset, input[1775:0] inp, output reg [221:0] outp); 

dsp_chain_4_int_sop_2_module inst_0 (.clk(clk),.reset(reset),.inp(inp[295:0]),.outp(outp[36:0])); 

dsp_chain_4_int_sop_2_module inst_1 (.clk(clk),.reset(reset),.inp(inp[591:296]),.outp(outp[73:37])); 

dsp_chain_4_int_sop_2_module inst_2 (.clk(clk),.reset(reset),.inp(inp[887:592]),.outp(outp[110:74])); 

dsp_chain_4_int_sop_2_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1183:888]),.outp(outp[147:111])); 

dsp_chain_4_int_sop_2_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1479:1184]),.outp(outp[184:148])); 

dsp_chain_4_int_sop_2_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1775:1480]),.outp(outp[221:185])); 

endmodule 

module fifo_256_40bit_module_24(input clk, input reset, input[1031:0] inp, output reg [1007:0] outp); 

fifo_256_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[42:0]),.outp(outp[41:0])); 

fifo_256_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[85:43]),.outp(outp[83:42])); 

fifo_256_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[128:86]),.outp(outp[125:84])); 

fifo_256_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[171:129]),.outp(outp[167:126])); 

fifo_256_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[214:172]),.outp(outp[209:168])); 

fifo_256_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[257:215]),.outp(outp[251:210])); 

fifo_256_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[300:258]),.outp(outp[293:252])); 

fifo_256_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[343:301]),.outp(outp[335:294])); 

fifo_256_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[386:344]),.outp(outp[377:336])); 

fifo_256_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[429:387]),.outp(outp[419:378])); 

fifo_256_40bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[472:430]),.outp(outp[461:420])); 

fifo_256_40bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[515:473]),.outp(outp[503:462])); 

fifo_256_40bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[558:516]),.outp(outp[545:504])); 

fifo_256_40bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[601:559]),.outp(outp[587:546])); 

fifo_256_40bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[644:602]),.outp(outp[629:588])); 

fifo_256_40bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[687:645]),.outp(outp[671:630])); 

fifo_256_40bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[730:688]),.outp(outp[713:672])); 

fifo_256_40bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[773:731]),.outp(outp[755:714])); 

fifo_256_40bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[816:774]),.outp(outp[797:756])); 

fifo_256_40bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[859:817]),.outp(outp[839:798])); 

fifo_256_40bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[902:860]),.outp(outp[881:840])); 

fifo_256_40bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[945:903]),.outp(outp[923:882])); 

fifo_256_40bit_module inst_22 (.clk(clk),.reset(reset),.inp(inp[988:946]),.outp(outp[965:924])); 

fifo_256_40bit_module inst_23 (.clk(clk),.reset(reset),.inp(inp[1031:989]),.outp(outp[1007:966])); 

endmodule 

module fifo_512_60bit_module_40(input clk, input reset, input[2519:0] inp, output reg [2479:0] outp); 

fifo_512_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[62:0]),.outp(outp[61:0])); 

fifo_512_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[125:63]),.outp(outp[123:62])); 

fifo_512_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[188:126]),.outp(outp[185:124])); 

fifo_512_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[251:189]),.outp(outp[247:186])); 

fifo_512_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[314:252]),.outp(outp[309:248])); 

fifo_512_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[377:315]),.outp(outp[371:310])); 

fifo_512_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[440:378]),.outp(outp[433:372])); 

fifo_512_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[503:441]),.outp(outp[495:434])); 

fifo_512_60bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[566:504]),.outp(outp[557:496])); 

fifo_512_60bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[629:567]),.outp(outp[619:558])); 

fifo_512_60bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[692:630]),.outp(outp[681:620])); 

fifo_512_60bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[755:693]),.outp(outp[743:682])); 

fifo_512_60bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[818:756]),.outp(outp[805:744])); 

fifo_512_60bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[881:819]),.outp(outp[867:806])); 

fifo_512_60bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[944:882]),.outp(outp[929:868])); 

fifo_512_60bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[1007:945]),.outp(outp[991:930])); 

fifo_512_60bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[1070:1008]),.outp(outp[1053:992])); 

fifo_512_60bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[1133:1071]),.outp(outp[1115:1054])); 

fifo_512_60bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[1196:1134]),.outp(outp[1177:1116])); 

fifo_512_60bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[1259:1197]),.outp(outp[1239:1178])); 

fifo_512_60bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[1322:1260]),.outp(outp[1301:1240])); 

fifo_512_60bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[1385:1323]),.outp(outp[1363:1302])); 

fifo_512_60bit_module inst_22 (.clk(clk),.reset(reset),.inp(inp[1448:1386]),.outp(outp[1425:1364])); 

fifo_512_60bit_module inst_23 (.clk(clk),.reset(reset),.inp(inp[1511:1449]),.outp(outp[1487:1426])); 

fifo_512_60bit_module inst_24 (.clk(clk),.reset(reset),.inp(inp[1574:1512]),.outp(outp[1549:1488])); 

fifo_512_60bit_module inst_25 (.clk(clk),.reset(reset),.inp(inp[1637:1575]),.outp(outp[1611:1550])); 

fifo_512_60bit_module inst_26 (.clk(clk),.reset(reset),.inp(inp[1700:1638]),.outp(outp[1673:1612])); 

fifo_512_60bit_module inst_27 (.clk(clk),.reset(reset),.inp(inp[1763:1701]),.outp(outp[1735:1674])); 

fifo_512_60bit_module inst_28 (.clk(clk),.reset(reset),.inp(inp[1826:1764]),.outp(outp[1797:1736])); 

fifo_512_60bit_module inst_29 (.clk(clk),.reset(reset),.inp(inp[1889:1827]),.outp(outp[1859:1798])); 

fifo_512_60bit_module inst_30 (.clk(clk),.reset(reset),.inp(inp[1952:1890]),.outp(outp[1921:1860])); 

fifo_512_60bit_module inst_31 (.clk(clk),.reset(reset),.inp(inp[2015:1953]),.outp(outp[1983:1922])); 

fifo_512_60bit_module inst_32 (.clk(clk),.reset(reset),.inp(inp[2078:2016]),.outp(outp[2045:1984])); 

fifo_512_60bit_module inst_33 (.clk(clk),.reset(reset),.inp(inp[2141:2079]),.outp(outp[2107:2046])); 

fifo_512_60bit_module inst_34 (.clk(clk),.reset(reset),.inp(inp[2204:2142]),.outp(outp[2169:2108])); 

fifo_512_60bit_module inst_35 (.clk(clk),.reset(reset),.inp(inp[2267:2205]),.outp(outp[2231:2170])); 

fifo_512_60bit_module inst_36 (.clk(clk),.reset(reset),.inp(inp[2330:2268]),.outp(outp[2293:2232])); 

fifo_512_60bit_module inst_37 (.clk(clk),.reset(reset),.inp(inp[2393:2331]),.outp(outp[2355:2294])); 

fifo_512_60bit_module inst_38 (.clk(clk),.reset(reset),.inp(inp[2456:2394]),.outp(outp[2417:2356])); 

fifo_512_60bit_module inst_39 (.clk(clk),.reset(reset),.inp(inp[2519:2457]),.outp(outp[2479:2418])); 

endmodule 

module fifo_256_60bit_module_18(input clk, input reset, input[1133:0] inp, output reg [1115:0] outp); 

fifo_256_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[62:0]),.outp(outp[61:0])); 

fifo_256_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[125:63]),.outp(outp[123:62])); 

fifo_256_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[188:126]),.outp(outp[185:124])); 

fifo_256_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[251:189]),.outp(outp[247:186])); 

fifo_256_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[314:252]),.outp(outp[309:248])); 

fifo_256_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[377:315]),.outp(outp[371:310])); 

fifo_256_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[440:378]),.outp(outp[433:372])); 

fifo_256_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[503:441]),.outp(outp[495:434])); 

fifo_256_60bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[566:504]),.outp(outp[557:496])); 

fifo_256_60bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[629:567]),.outp(outp[619:558])); 

fifo_256_60bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[692:630]),.outp(outp[681:620])); 

fifo_256_60bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[755:693]),.outp(outp[743:682])); 

fifo_256_60bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[818:756]),.outp(outp[805:744])); 

fifo_256_60bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[881:819]),.outp(outp[867:806])); 

fifo_256_60bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[944:882]),.outp(outp[929:868])); 

fifo_256_60bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[1007:945]),.outp(outp[991:930])); 

fifo_256_60bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[1070:1008]),.outp(outp[1053:992])); 

fifo_256_60bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[1133:1071]),.outp(outp[1115:1054])); 

endmodule 

module fifo_512_40bit_module_26(input clk, input reset, input[1117:0] inp, output reg [1091:0] outp); 

fifo_512_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[42:0]),.outp(outp[41:0])); 

fifo_512_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[85:43]),.outp(outp[83:42])); 

fifo_512_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[128:86]),.outp(outp[125:84])); 

fifo_512_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[171:129]),.outp(outp[167:126])); 

fifo_512_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[214:172]),.outp(outp[209:168])); 

fifo_512_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[257:215]),.outp(outp[251:210])); 

fifo_512_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[300:258]),.outp(outp[293:252])); 

fifo_512_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[343:301]),.outp(outp[335:294])); 

fifo_512_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[386:344]),.outp(outp[377:336])); 

fifo_512_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[429:387]),.outp(outp[419:378])); 

fifo_512_40bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[472:430]),.outp(outp[461:420])); 

fifo_512_40bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[515:473]),.outp(outp[503:462])); 

fifo_512_40bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[558:516]),.outp(outp[545:504])); 

fifo_512_40bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[601:559]),.outp(outp[587:546])); 

fifo_512_40bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[644:602]),.outp(outp[629:588])); 

fifo_512_40bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[687:645]),.outp(outp[671:630])); 

fifo_512_40bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[730:688]),.outp(outp[713:672])); 

fifo_512_40bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[773:731]),.outp(outp[755:714])); 

fifo_512_40bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[816:774]),.outp(outp[797:756])); 

fifo_512_40bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[859:817]),.outp(outp[839:798])); 

fifo_512_40bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[902:860]),.outp(outp[881:840])); 

fifo_512_40bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[945:903]),.outp(outp[923:882])); 

fifo_512_40bit_module inst_22 (.clk(clk),.reset(reset),.inp(inp[988:946]),.outp(outp[965:924])); 

fifo_512_40bit_module inst_23 (.clk(clk),.reset(reset),.inp(inp[1031:989]),.outp(outp[1007:966])); 

fifo_512_40bit_module inst_24 (.clk(clk),.reset(reset),.inp(inp[1074:1032]),.outp(outp[1049:1008])); 

fifo_512_40bit_module inst_25 (.clk(clk),.reset(reset),.inp(inp[1117:1075]),.outp(outp[1091:1050])); 

endmodule 

module dsp_chain_3_int_sop_2_module_16(input clk, input reset, input[3551:0] inp, output reg [591:0] outp); 

dsp_chain_3_int_sop_2_module inst_0 (.clk(clk),.reset(reset),.inp(inp[221:0]),.outp(outp[36:0])); 

dsp_chain_3_int_sop_2_module inst_1 (.clk(clk),.reset(reset),.inp(inp[443:222]),.outp(outp[73:37])); 

dsp_chain_3_int_sop_2_module inst_2 (.clk(clk),.reset(reset),.inp(inp[665:444]),.outp(outp[110:74])); 

dsp_chain_3_int_sop_2_module inst_3 (.clk(clk),.reset(reset),.inp(inp[887:666]),.outp(outp[147:111])); 

dsp_chain_3_int_sop_2_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1109:888]),.outp(outp[184:148])); 

dsp_chain_3_int_sop_2_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1331:1110]),.outp(outp[221:185])); 

dsp_chain_3_int_sop_2_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1553:1332]),.outp(outp[258:222])); 

dsp_chain_3_int_sop_2_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1775:1554]),.outp(outp[295:259])); 

dsp_chain_3_int_sop_2_module inst_8 (.clk(clk),.reset(reset),.inp(inp[1997:1776]),.outp(outp[332:296])); 

dsp_chain_3_int_sop_2_module inst_9 (.clk(clk),.reset(reset),.inp(inp[2219:1998]),.outp(outp[369:333])); 

dsp_chain_3_int_sop_2_module inst_10 (.clk(clk),.reset(reset),.inp(inp[2441:2220]),.outp(outp[406:370])); 

dsp_chain_3_int_sop_2_module inst_11 (.clk(clk),.reset(reset),.inp(inp[2663:2442]),.outp(outp[443:407])); 

dsp_chain_3_int_sop_2_module inst_12 (.clk(clk),.reset(reset),.inp(inp[2885:2664]),.outp(outp[480:444])); 

dsp_chain_3_int_sop_2_module inst_13 (.clk(clk),.reset(reset),.inp(inp[3107:2886]),.outp(outp[517:481])); 

dsp_chain_3_int_sop_2_module inst_14 (.clk(clk),.reset(reset),.inp(inp[3329:3108]),.outp(outp[554:518])); 

dsp_chain_3_int_sop_2_module inst_15 (.clk(clk),.reset(reset),.inp(inp[3551:3330]),.outp(outp[591:555])); 

endmodule 


module fifo_256_40bit_module_4(input clk, input reset, input[171:0] inp, output reg [167:0] outp); 

fifo_256_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[42:0]),.outp(outp[41:0])); 

fifo_256_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[85:43]),.outp(outp[83:42])); 

fifo_256_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[128:86]),.outp(outp[125:84])); 

fifo_256_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[171:129]),.outp(outp[167:126])); 

endmodule 

module dsp_chain_4_int_sop_2_module_8(input clk, input reset, input[2367:0] inp, output reg [295:0] outp); 

dsp_chain_4_int_sop_2_module inst_0 (.clk(clk),.reset(reset),.inp(inp[295:0]),.outp(outp[36:0])); 

dsp_chain_4_int_sop_2_module inst_1 (.clk(clk),.reset(reset),.inp(inp[591:296]),.outp(outp[73:37])); 

dsp_chain_4_int_sop_2_module inst_2 (.clk(clk),.reset(reset),.inp(inp[887:592]),.outp(outp[110:74])); 

dsp_chain_4_int_sop_2_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1183:888]),.outp(outp[147:111])); 

dsp_chain_4_int_sop_2_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1479:1184]),.outp(outp[184:148])); 

dsp_chain_4_int_sop_2_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1775:1480]),.outp(outp[221:185])); 

dsp_chain_4_int_sop_2_module inst_6 (.clk(clk),.reset(reset),.inp(inp[2071:1776]),.outp(outp[258:222])); 

dsp_chain_4_int_sop_2_module inst_7 (.clk(clk),.reset(reset),.inp(inp[2367:2072]),.outp(outp[295:259])); 

endmodule 

module tensor_block_int8_module_1(input clk, input reset, input[264:0] inp, output reg [250:0] outp); 

tensor_block_int8_module inst_0 (.clk(clk),.reset(reset),.inp(inp[264:0]),.outp(outp[250:0])); 

endmodule 

module fifo_512_60bit_module_32(input clk, input reset, input[2015:0] inp, output reg [1983:0] outp); 

fifo_512_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[62:0]),.outp(outp[61:0])); 

fifo_512_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[125:63]),.outp(outp[123:62])); 

fifo_512_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[188:126]),.outp(outp[185:124])); 

fifo_512_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[251:189]),.outp(outp[247:186])); 

fifo_512_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[314:252]),.outp(outp[309:248])); 

fifo_512_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[377:315]),.outp(outp[371:310])); 

fifo_512_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[440:378]),.outp(outp[433:372])); 

fifo_512_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[503:441]),.outp(outp[495:434])); 

fifo_512_60bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[566:504]),.outp(outp[557:496])); 

fifo_512_60bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[629:567]),.outp(outp[619:558])); 

fifo_512_60bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[692:630]),.outp(outp[681:620])); 

fifo_512_60bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[755:693]),.outp(outp[743:682])); 

fifo_512_60bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[818:756]),.outp(outp[805:744])); 

fifo_512_60bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[881:819]),.outp(outp[867:806])); 

fifo_512_60bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[944:882]),.outp(outp[929:868])); 

fifo_512_60bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[1007:945]),.outp(outp[991:930])); 

fifo_512_60bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[1070:1008]),.outp(outp[1053:992])); 

fifo_512_60bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[1133:1071]),.outp(outp[1115:1054])); 

fifo_512_60bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[1196:1134]),.outp(outp[1177:1116])); 

fifo_512_60bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[1259:1197]),.outp(outp[1239:1178])); 

fifo_512_60bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[1322:1260]),.outp(outp[1301:1240])); 

fifo_512_60bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[1385:1323]),.outp(outp[1363:1302])); 

fifo_512_60bit_module inst_22 (.clk(clk),.reset(reset),.inp(inp[1448:1386]),.outp(outp[1425:1364])); 

fifo_512_60bit_module inst_23 (.clk(clk),.reset(reset),.inp(inp[1511:1449]),.outp(outp[1487:1426])); 

fifo_512_60bit_module inst_24 (.clk(clk),.reset(reset),.inp(inp[1574:1512]),.outp(outp[1549:1488])); 

fifo_512_60bit_module inst_25 (.clk(clk),.reset(reset),.inp(inp[1637:1575]),.outp(outp[1611:1550])); 

fifo_512_60bit_module inst_26 (.clk(clk),.reset(reset),.inp(inp[1700:1638]),.outp(outp[1673:1612])); 

fifo_512_60bit_module inst_27 (.clk(clk),.reset(reset),.inp(inp[1763:1701]),.outp(outp[1735:1674])); 

fifo_512_60bit_module inst_28 (.clk(clk),.reset(reset),.inp(inp[1826:1764]),.outp(outp[1797:1736])); 

fifo_512_60bit_module inst_29 (.clk(clk),.reset(reset),.inp(inp[1889:1827]),.outp(outp[1859:1798])); 

fifo_512_60bit_module inst_30 (.clk(clk),.reset(reset),.inp(inp[1952:1890]),.outp(outp[1921:1860])); 

fifo_512_60bit_module inst_31 (.clk(clk),.reset(reset),.inp(inp[2015:1953]),.outp(outp[1983:1922])); 

endmodule 

module dsp_chain_2_int_sop_2_module_25(input clk, input reset, input[3699:0] inp, output reg [924:0] outp); 

dsp_chain_2_int_sop_2_module inst_0 (.clk(clk),.reset(reset),.inp(inp[147:0]),.outp(outp[36:0])); 

dsp_chain_2_int_sop_2_module inst_1 (.clk(clk),.reset(reset),.inp(inp[295:148]),.outp(outp[73:37])); 

dsp_chain_2_int_sop_2_module inst_2 (.clk(clk),.reset(reset),.inp(inp[443:296]),.outp(outp[110:74])); 

dsp_chain_2_int_sop_2_module inst_3 (.clk(clk),.reset(reset),.inp(inp[591:444]),.outp(outp[147:111])); 

dsp_chain_2_int_sop_2_module inst_4 (.clk(clk),.reset(reset),.inp(inp[739:592]),.outp(outp[184:148])); 

dsp_chain_2_int_sop_2_module inst_5 (.clk(clk),.reset(reset),.inp(inp[887:740]),.outp(outp[221:185])); 

dsp_chain_2_int_sop_2_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1035:888]),.outp(outp[258:222])); 

dsp_chain_2_int_sop_2_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1183:1036]),.outp(outp[295:259])); 

dsp_chain_2_int_sop_2_module inst_8 (.clk(clk),.reset(reset),.inp(inp[1331:1184]),.outp(outp[332:296])); 

dsp_chain_2_int_sop_2_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1479:1332]),.outp(outp[369:333])); 

dsp_chain_2_int_sop_2_module inst_10 (.clk(clk),.reset(reset),.inp(inp[1627:1480]),.outp(outp[406:370])); 

dsp_chain_2_int_sop_2_module inst_11 (.clk(clk),.reset(reset),.inp(inp[1775:1628]),.outp(outp[443:407])); 

dsp_chain_2_int_sop_2_module inst_12 (.clk(clk),.reset(reset),.inp(inp[1923:1776]),.outp(outp[480:444])); 

dsp_chain_2_int_sop_2_module inst_13 (.clk(clk),.reset(reset),.inp(inp[2071:1924]),.outp(outp[517:481])); 

dsp_chain_2_int_sop_2_module inst_14 (.clk(clk),.reset(reset),.inp(inp[2219:2072]),.outp(outp[554:518])); 

dsp_chain_2_int_sop_2_module inst_15 (.clk(clk),.reset(reset),.inp(inp[2367:2220]),.outp(outp[591:555])); 

dsp_chain_2_int_sop_2_module inst_16 (.clk(clk),.reset(reset),.inp(inp[2515:2368]),.outp(outp[628:592])); 

dsp_chain_2_int_sop_2_module inst_17 (.clk(clk),.reset(reset),.inp(inp[2663:2516]),.outp(outp[665:629])); 

dsp_chain_2_int_sop_2_module inst_18 (.clk(clk),.reset(reset),.inp(inp[2811:2664]),.outp(outp[702:666])); 

dsp_chain_2_int_sop_2_module inst_19 (.clk(clk),.reset(reset),.inp(inp[2959:2812]),.outp(outp[739:703])); 

dsp_chain_2_int_sop_2_module inst_20 (.clk(clk),.reset(reset),.inp(inp[3107:2960]),.outp(outp[776:740])); 

dsp_chain_2_int_sop_2_module inst_21 (.clk(clk),.reset(reset),.inp(inp[3255:3108]),.outp(outp[813:777])); 

dsp_chain_2_int_sop_2_module inst_22 (.clk(clk),.reset(reset),.inp(inp[3403:3256]),.outp(outp[850:814])); 

dsp_chain_2_int_sop_2_module inst_23 (.clk(clk),.reset(reset),.inp(inp[3551:3404]),.outp(outp[887:851])); 

dsp_chain_2_int_sop_2_module inst_24 (.clk(clk),.reset(reset),.inp(inp[3699:3552]),.outp(outp[924:888])); 

endmodule 

module fifo_256_40bit_module_6(input clk, input reset, input[257:0] inp, output reg [251:0] outp); 

fifo_256_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[42:0]),.outp(outp[41:0])); 

fifo_256_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[85:43]),.outp(outp[83:42])); 

fifo_256_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[128:86]),.outp(outp[125:84])); 

fifo_256_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[171:129]),.outp(outp[167:126])); 

fifo_256_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[214:172]),.outp(outp[209:168])); 

fifo_256_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[257:215]),.outp(outp[251:210])); 

endmodule 
module adder_tree_1_16bit (input clk,input reset,input [31:0] inp, output reg [31:0] outp);

adder_tree_1stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.sum_out(outp));

endmodule

module adder_tree_2_16bit (input clk, input reset, input [63:0] inp, output reg [31:0] outp);

adder_tree_2stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.sum_out(outp));

endmodule

module adder_tree_3_16bit (input clk, input reset, input [127:0] inp, output reg [31:0] outp);

adder_tree_3stage_16bit inst (.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.inp20(inp[79:64]),.inp21(inp[95:80]),.inp30(inp[111:96]),.inp31(inp[127:112]),.sum_out(outp));

endmodule

module adder_tree_4_16bit (input clk, input reset, input [255:0] inp, output reg [31:0] outp);

adder_tree_4stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.inp20(inp[79:64]),.inp21(inp[95:80]),.inp30(inp[111:96]),.inp31(inp[127:112]),.inp40(inp[143:128]),.inp41(inp[159:144]),.inp50(inp[175:160]),.inp51(inp[191:176]),.inp60(inp[207:192]),.inp61(inp[223:208]),.inp70(inp[239:224]),.inp71(inp[255:240]),.sum_out(outp));

endmodule

module adder_tree_1_8bit (input clk, input reset, input [15:0] inp, output reg [15:0] outp);

adder_tree_1stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.sum_out(outp));

endmodule

module adder_tree_2_8bit (input clk, input reset, input [31:0] inp, output reg [15:0] outp);

adder_tree_2stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.sum_out(outp));

endmodule

module adder_tree_3_8bit (input clk, input reset, input [63:0] inp, output reg [15:0] outp);

adder_tree_3stage_8bit inst (.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.inp20(inp[39:32]),.inp21(inp[47:40]),.inp30(inp[55:48]),.inp31(inp[63:56]),.sum_out(outp));

endmodule

module adder_tree_4_8bit (input clk, input reset, input [127:0] inp, output reg [15:0] outp);

adder_tree_4stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.inp20(inp[39:32]),.inp21(inp[47:40]),.inp30(inp[55:48]),.inp31(inp[63:56]),.inp40(inp[71:64]),.inp41(inp[79:72]),.inp50(inp[87:80]),.inp51(inp[95:88]),.inp60(inp[103:96]),.inp61(inp[111:104]),.inp70(inp[119:112]),.inp71(inp[127:120]),.sum_out(outp));

endmodule

module adder_tree_1_4bit (input clk, input reset, input [7:0] inp, output reg [7:0] outp);

adder_tree_1stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.sum_out(outp));

endmodule

module adder_tree_2_4bit (input clk, input reset, input [15:0] inp, output reg [7:0] outp);

adder_tree_2stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.sum_out(outp));

endmodule

module adder_tree_3_4bit (input clk, input reset, input [31:0] inp, output reg [7:0] outp);

adder_tree_3stage_4bit inst (.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.inp20(inp[19:16]),.inp21(inp[23:20]),.inp30(inp[27:24]),.inp31(inp[31:28]),.sum_out(outp));

endmodule

module adder_tree_4_4bit (input clk, input reset, input [63:0] inp, output reg [7:0] outp);

adder_tree_4stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.inp20(inp[19:16]),.inp21(inp[23:20]),.inp30(inp[27:24]),.inp31(inp[31:28]),.inp40(inp[35:32]),.inp41(inp[39:36]),.inp50(inp[43:40]),.inp51(inp[47:44]),.inp60(inp[51:48]),.inp61(inp[55:52]),.inp70(inp[59:56]),.inp71(inp[63:60]),.sum_out(outp));

endmodule

module adder_tree_3_fp16bit (input clk, input reset, input [131:0] inp, output reg [15:0] outp);

mode4_adder_tree inst(
  .inp0(inp[15:0]),
  .inp1(inp[31:16]),
  .inp2(inp[47:32]),
  .inp3(inp[63:48]),
  .inp4(inp[79:64]),
  .inp5(inp[95:80]),
  .inp6(inp[111:96]),
  .inp7(inp[127:112]),
  .mode4_stage0_run(inp[128]),
  .mode4_stage1_run(inp[129]),
  .mode4_stage2_run(inp[130]),
  .mode4_stage3_run(inp[131]),

  .clk(clk),
  .reset(reset),
  .outp(outp[15:0])
);

endmodule

module dpram_1024_32bit_module (input clk, input reset, input [85:0] inp, output reg [63:0] outp);

dpram inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[53:22]),.data_b(inp[85:54]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_1024_64bit_module (input clk, input reset, input [149:0] inp, output reg [63:0] outp );

dpram_1024_64bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[85:22]),.data_b(inp[149:86]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_2048_64bit_module (input clk, input reset, input [151:0] inp, output reg [127:0] outp);

dpram_2048_64bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[87:24]),.data_b(inp[151:88]),.out_a(outp[63:0]),.out_b(outp[127:64]));

endmodule

module dpram_2048_32bit_module (input clk, input reset, input [87:0] inp, output reg [63:0] outp);

dpram_2048_32bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[55:24]),.data_b(inp[87:56]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_1024_40bit_module (input clk, input reset, input [101:0] inp, output reg [79:0] outp);

dpram_1024_40bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[61:22]),.data_b(inp[101:62]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_1024_60bit_module (input clk, input reset, input [141:0] inp, output reg [119:0] outp);

dpram_1024_60bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[81:22]),.data_b(inp[141:82]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dpram_2048_40bit_module (input clk, input reset, input [103:0] inp, output reg [79:0] outp);

dpram_2048_40bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[63:24]),.data_b(inp[103:64]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_2048_60bit_module (input clk, input reset, input [143:0] inp, output reg [119:0] outp);

dpram_2048_60bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[83:24]),.data_b(inp[143:84]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dpram_4096_40bit_module (input clk, input reset, input [105:0] inp, output reg [79:0] outp);

dpram_4096_40bit inst (.clk(clk),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[65:26]),.data_b(inp[105:66]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_4096_60bit_module (input clk, input reset, input [145:0] inp, output reg [119:0] outp);

dpram_4096_60bit inst (.clk(clk),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[85:26]),.data_b(inp[145:86]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module spram_1024_32bit_module (input clk,input reset,input [42:0] inp, output reg [31:0] outp);

spram inst (.clk(clk),.address(inp[9:0]),.wren(inp[10]),.data(inp[42:11]),.out(outp));

endmodule

module spram_2048_40bit_module (input clk,input reset,input [51:0] inp, output reg [39:0] outp);

spram_2048_40bit inst (.clk(clk),.address(inp[10:0]),.wren(inp[11]),.data(inp[51:12]),.out(outp));

endmodule

module spram_2048_60bit_module (input clk,input reset,input [71:0] inp, output reg [59:0] outp);

spram_2048_60bit inst (.clk(clk),.address(inp[10:0]),.wren(inp[11]),.data(inp[71:12]),.out(outp));

endmodule

module spram_4096_40bit_module (input clk,input reset,input [52:0] inp, output reg [39:0] outp);

spram_4096_40bit inst (.clk(clk),.address(inp[11:0]),.wren(inp[12]),.data(inp[52:13]),.out(outp));

endmodule

module spram_4096_60bit_module (input clk,input reset,input [72:0] inp, output reg [59:0] outp);

spram_4096_60bit inst (.clk(clk),.address(inp[11:0]),.wren(inp[12]),.data(inp[72:13]),.out(outp));

endmodule

module dbram_2048_40bit_module (input clk,input reset,input [103:0] inp, output reg [79:0] outp);

dbram_2048_40bit inst (.clk(clk),.reset(reset),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[63:24]),.data_b(inp[103:64]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dbram_2048_60bit_module (input clk,input reset,input [143:0] inp, output reg [119:0] outp);

dbram_2048_60bit inst (.clk(clk),.reset(reset),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[83:24]),.data_b(inp[143:84]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dbram_4096_40bit_module (input clk,input reset,input [105:0] inp, output reg [79:0] outp);

dbram_4096_40bit inst (.clk(clk),.reset(reset),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[65:26]),.data_b(inp[105:66]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dbram_4096_60bit_module (input clk,input reset,input [145:0] inp, output reg [119:0] outp);

dbram_4096_60bit inst (.clk(clk),.reset(reset),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[85:26]),.data_b(inp[145:86]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule


module fifo_256_40bit_module (input clk,input reset,input [42:0] inp, output reg [41:0] outp);

fifo_256_40bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[40:1]),.we(inp[41]),.dout(outp[39:0]),.re(inp[42]),.full(outp[40]),.empty(outp[41]));

endmodule

module fifo_256_60bit_module (input clk,input reset,input [62:0] inp, output reg [61:0] outp);

fifo_256_60bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[60:1]),.we(inp[61]),.dout(outp[59:0]),.re(inp[62]),.full(outp[60]),.empty(outp[61]));

endmodule

module fifo_512_60bit_module (input clk,input reset,input [62:0] inp, output reg [61:0] outp);

fifo_512_60bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[60:1]),.we(inp[61]),.dout(outp[59:0]),.re(inp[62]),.full(outp[60]),.empty(outp[61]));

endmodule

module fifo_512_40bit_module (input clk,input reset,input [42:0] inp, output reg [41:0] outp);

fifo_512_40bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[40:1]),.we(inp[41]),.dout(outp[39:0]),.re(inp[42]),.full(outp[40]),.empty(outp[41]));

endmodule

module tanh_16bit (input clk,input reset, input [15:0] inp, output reg [15:0] outp);

tanh inst (.x(inp),.tanh_out(outp));

endmodule

module sigmoid_16bit (input clk,input reset, input [15:0] inp, output reg [15:0] outp);

sigmoid inst (.x(inp),.sig_out(outp));

endmodule

module systolic_array_4_16bit (input clk, input reset, input [254:0] inp, output reg [130:0] outp);

matmul_4x4_systolic inst(
 .clk(clk),
 .reset(inp[254]),
 .pe_reset(reset),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[11:1]),
 .address_mat_b(inp[22:12]),
 .address_mat_c(inp[33:23]),
 .address_stride_a(inp[41:34]),
 .address_stride_b(inp[49:42]),
 .address_stride_c(inp[57:50]),
 .a_data(inp[89:58]),
 .b_data(inp[121:90]),
 .a_data_in(inp[153:122]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[185:154]),
 .c_data_in(inp[217:186]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[32:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[64:33]),
 .b_data_out(outp[96:65]),
 .a_addr(outp[107:97]),
 .b_addr(outp[118:108]),
 .c_addr(outp[129:119]),
 .c_data_available(outp[130]),
 .validity_mask_a_rows(inp[221:218]),
 .validity_mask_a_cols_b_rows(inp[225:222]),
 .validity_mask_b_cols(inp[229:226]),
 .final_mat_mul_size(inp[237:230]),
 .a_loc(inp[245:238]),
 .b_loc(inp[253:246])
);

endmodule

module systolic_array_8_16bit (input clk, input reset, input [785:0] inp, output reg [433:0] outp);

matmul_8x8_systolic inst(
 .clk(clk),
 .reset(reset),
 .pe_reset(inp[785]),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[16:1]),
 .address_mat_b(inp[32:17]),
 .address_mat_c(inp[48:33]),
 .address_stride_a(inp[64:49]),
 .address_stride_b(inp[80:65]),
 .address_stride_c(inp[96:81]),
 .a_data(inp[224:97]),
 .b_data(inp[352:225]),
 .a_data_in(inp[480:353]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[608:481]),
 .c_data_in(inp[736:609]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[128:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[256:129]),
 .b_data_out(outp[384:257]),
 .a_addr(outp[400:385]),
 .b_addr(outp[416:401]),
 .c_addr(outp[432:417]),
 .c_data_available(outp[433]),
 .validity_mask_a_rows(inp[744:737]),
 .validity_mask_a_cols_b_rows(inp[752:745]),
 .validity_mask_b_cols(inp[760:753]),
 .final_mat_mul_size(inp[768:761]),
 .a_loc(inp[776:769]),
 .b_loc(inp[784:777])
);

endmodule

module systolic_array_4_fp16bit (input clk, input reset, input [417:0] inp, output reg [223:0] outp);

matmul_4x4_fp_systolic inst(
 .clk(clk),
 .reset(reset),
 .pe_reset(inp[417]),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[10:1]),
 .address_mat_b(inp[20:11]),
 .address_mat_c(inp[30:21]),
 .address_stride_a(inp[40:31]),
 .address_stride_b(inp[50:41]),
 .address_stride_c(inp[60:51]),
 .a_data(inp[124:61]),
 .b_data(inp[188:125]),
 .a_data_in(inp[252:189]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[316:253]),
 .c_data_in(inp[380:317]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[64:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[128:65]),
 .b_data_out(outp[192:129]),
 .a_addr(outp[202:193]),
 .b_addr(outp[212:203]),
 .c_addr(outp[222:213]),
 .c_data_available(outp[223]),
 .validity_mask_a_rows(inp[384:381]),
 .validity_mask_a_cols_b_rows(inp[388:385]),
 .validity_mask_b_cols(inp[392:389]),
 .final_mat_mul_size(inp[400:393]),
 .a_loc(inp[408:401]),
 .b_loc(inp[416:409])
);

endmodule

module dsp_chain_2_int_sop_2_module (input clk, input reset, input [147:0] inp, output reg [36:0] outp);

dsp_chain_2_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.result(outp[36:0]));

endmodule

module dsp_chain_3_int_sop_2_module (input clk, input reset, input [221:0] inp, output reg [36:0] outp);

dsp_chain_3_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.ax3(inp[165:148]),.ay3(inp[184:166]),.bx3(inp[202:185]),.by3(inp[221:203]),.result(outp[36:0]));

endmodule

module dsp_chain_4_int_sop_2_module (input clk, input reset, input [295:0] inp, output reg [36:0] outp);

dsp_chain_4_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.ax3(inp[165:148]),.ay3(inp[184:166]),.bx3(inp[202:185]),.by3(inp[221:203]),.ax4(inp[239:222]),.ay4(inp[258:240]),.bx4(inp[276:259]),.by4(inp[295:277]),.result(outp[36:0]));

endmodule

module dsp_chain_2_fp16_sop2_mult_module (input clk, input reset, input [127:0] inp, output reg [31:0] outp);

dsp_chain_2_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.result(outp));

endmodule

module dsp_chain_3_fp16_sop2_mult_module (input clk, input reset, input [191:0] inp, output reg [31:0] outp);

dsp_chain_3_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.top_a3(inp[143:128]),.top_b3(inp[159:144]),.bot_a3(inp[175:160]),.bot_b3(inp[191:176]),.result(outp));

endmodule

module dsp_chain_4_fp16_sop2_mult_module (input clk, input reset, input [255:0] inp, output reg [31:0] outp);

dsp_chain_4_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.top_a3(inp[143:128]),.top_b3(inp[159:144]),.bot_a3(inp[175:160]),.bot_b3(inp[191:176]),.top_a4(inp[207:192]),.top_b4(inp[223:208]),.bot_a4(inp[239:224]),.bot_b4(inp[255:240]),.result(outp));

endmodule

module tensor_block_bf16_module (input clk, input reset, input [264:0] inp, output reg [271:0] outp);

tensor_block_bf16 inst(
	.clk(clk),
	.reset(reset),

	.data_in(inp[79:0]),
	.cascade_in(inp[159:80]),
	.acc0_in(inp[191:160]),
	.acc1_in(inp[223:192]),
	.acc2_in(inp[255:224]),
	.accumulator_input1_select(inp[258:256]),

	.out0(outp[31:0]),
	.out1(outp[63:32]),
	.out2(outp[95:64]),
	.cascade_out(outp[175:96]),
	.acc0_out(outp[207:176]),
	.acc1_out(outp[239:208]),
	.acc2_out(outp[271:240]),

	.mux1_select(inp[259]),
	.dot_unit_input_1_enable(inp[260]),
	.bank0_data_in_enable(inp[261]),
	.bank1_data_in_enable(inp[262]),
	.cascade_out_select(inp[263]),
	.dot_unit_input_2_select(inp[264])

	);

endmodule

module tensor_block_int8_module (input clk, input reset, input [264:0] inp, output reg [250:0] outp);

tensor_block inst(
	.clk(clk),
	.reset(reset),

	.data_in(inp[79:0]),
	.cascade_in(inp[159:80]),
	.acc0_in(inp[191:160]),
	.acc1_in(inp[223:192]),
	.acc2_in(inp[255:224]),
	.accumulator_input1_select(inp[258:256]),

	.out0(outp[24:0]),
	.out1(outp[49:25]),
	.out2(outp[74:50]),
	.cascade_out(outp[154:75]),
	.acc0_out(outp[186:155]),
	.acc1_out(outp[218:187]),
	.acc2_out(outp[250:219]),

	.mux1_select(inp[259]),
	.dot_unit_input_1_enable(inp[260]),
	.bank0_data_in_enable(inp[261]),
	.bank1_data_in_enable(inp[262]),
	.cascade_out_select(inp[263]),
	.dot_unit_input_2_select(inp[264])

	);

endmodule


module activation_32_8bit_module (input clk, input reset, input [260:0] inp, output reg [257:0] outp);

activation_32_8bit inst (
    .activation_type(inp[0]),
    .enable_activation(inp[1]),
    .in_data_available(inp[2]),
    .inp_data(inp[258:3]),
    .out_data(outp[255:0]),
    .out_data_available(outp[256]),
    .validity_mask(inp[260:259]),
    .done_activation(outp[257]),
    .clk(clk),
    .reset(reset)
);

endmodule

module activation_32_16bit_module (input clk, input reset, input [515:0] inp, output reg [513:0] outp);

activation_32_16bit inst (
    .activation_type(inp[0]),
    .enable_activation(inp[1]),
    .in_data_available(inp[2]),
    .inp_data(inp[514:3]),
    .out_data(outp[511:0]),
    .out_data_available(outp[512]),
    .validity_mask(inp[515:514]),
    .done_activation(outp[513]),
    .clk(clk),
    .reset(reset)
);

endmodule

module fsm(input clk, input reset, input i1, input i2, output reg o);
// mealy machine

reg [1:0] current_state; 
reg [1:0] next_state;

wire [1:0] inp; 
assign inp = {i2,i1}; 

always@(posedge clk) begin 
	if (reset == 1'b1) begin 
		current_state <= 1'b0; 
	end
	else begin 
		current_state <= next_state; 
	end
end

always@(posedge clk) begin 

	next_state = current_state; 

	case(current_state)
		2'b00:	begin 
							if(inp == 2'b00) begin 
								next_state <= 2'b00; 
								o <= 1'b0; 
							end
							if (inp == 2'b01) begin 
								next_state <= 2'b11;
								o <= 1'b1;
							end
							if(inp == 2'b10) begin
  							next_state <= 2'b01;
  							o <= 1'b0;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b10;
							  o <= 1'b0;
							end
					 	end 
		2'b01:	begin 
							if(inp == 2'b00) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b01;
							  o <= 1'b0;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b00;
							  o <= 1'b1;
							end
						end
		2'b10:	begin 
							if(inp == 2'b00) begin
							  next_state <= 2'b11;
							  o <= 1'b0;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b11;
							  o <= 1'b0;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
						end
		2'b11:	begin 
							if(inp == 2'b00) begin
  							next_state <= 2'b00;
							  o <= 1'b1;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b11;
							  o <= 1'b1;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
						end
//		defualt:	begin  
//								next_state <= 2'b00;
//								o <= 1'b0; 
//							end
	endcase
end 

endmodule 
module xor_module (input clk, input reset, input i1, input i2, output reg o);

always@(posedge clk) begin 
if (reset ==1'b1) begin 
o<= 1'b0; 
end
else begin
o <= i1^i2; 
end 
end
endmodule
module mux_module (input clk, input reset, input i1, input i2, output reg o, input sel);

always@(posedge clk) begin 
if (reset ==1'b1) begin 
	o<= 1'b0; 
end

else begin
	if (sel == 1'b0) begin 
		o <= i1;
	end
	else begin
		o <= i2; 
	end 
end 

end

endmodule

`ifdef complex_dsp
module int_sop_2_dspchain (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
	chainin,
	resulta,
	chainout);
input [10:0] mode_sigs;
input clk;
input reset; 
input [17:0] ax, bx;
input [18:0] ay, by;
input [36:0] chainin;

output reg [36:0] resulta;
output reg [36:0] chainout;

wire [11:0] mode_sigs_int;
assign mode_sigs_int = {1'b0, mode_sigs};

int_sop_2 inst1(.clk(clk),.reset(reset),.ax(ax),.bx(bx),.ay(ay),.by(by),.mode_sigs(mode_sigs_int),.chainin(chainin),.result(resulta),.chainout(chainout)); 

endmodule
`else
module int_sop_2_dspchain (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
	chainin,
	resulta,
	chainout);
input [10:0] mode_sigs;
input clk;
input reset; 
input [17:0] ax, bx;
input [18:0] ay, by;
input [36:0] chainin;

output reg [36:0] resulta;
output reg [36:0] chainout;
reg [17:0] ax_reg;
reg [18:0] ay_reg;
reg [17:0] bx_reg;
reg [18:0] by_reg;
reg [36:0] resulta;
always @(posedge clk) begin
  if(reset) begin
    resulta <= 0;
    ax_reg <= 0;
    ay_reg <= 0;
    bx_reg <= 0;
    by_reg <= 0;
  end
  else begin
    ax_reg <= ax;
    ay_reg <= ay;
    bx_reg <= bx;
    by_reg <= by;
    resulta <= ax_reg * ay_reg + bx_reg * by_reg + chainin;
  end
end
assign chainout = resulta;
endmodule
`endif

`ifdef complex_dsp
module fp16_sop2_mult_dspchain (clk,reset,top_a,top_b,bot_a,bot_b,fp32_in,mode_sigs,chainin,chainout,result);
input clk; 
input reset;
input [10:0] mode_sigs; 
input [15:0] top_a,top_b,bot_a,bot_b;
input [31:0] chainin,fp32_in; 
output reg [31:0] chainout, result;

fp16_sop2_mult inst1(.clk(clk),.reset(reset),.top_a(top_a),.top_b(top_b),.bot_a(bot_a),.bot_b(bot_b),.fp32_in(fp32_in),.mode_sigs(mode_sigs),.chainin(chainin),.chainout(chainout),.result(result)); 

endmodule

`else
module fp16_sop2_mult_dspchain (clk,reset,top_a,top_b,bot_a,bot_b,fp32_in,mode_sigs,chainin,chainout,result);
input clk; 
input reset;
input [10:0] mode_sigs; 
input [15:0] top_a,top_b,bot_a,bot_b;
input [31:0] chainin,fp32_in; 
output reg [31:0] chainout, result; 

reg [15:0] top_a_reg,top_b_reg,bot_a_reg,bot_b_reg; 
reg [31:0] chainin_reg; 
reg [31:0] r1,r2,r3; 
always@(posedge clk) begin 
if(reset) begin 
top_a_reg<= 16'b0; 
top_b_reg<= 16'b0; 
bot_a_reg<= 16'b0; 
bot_b_reg<= 16'b0;
//result<=32'b0;
//chainout<=32'b0;
chainin_reg<=32'b0;   
end
else begin 
top_a_reg<=top_a; 
top_b_reg<=top_b; 
bot_a_reg<=bot_a;
bot_b_reg<=bot_b;
//chainout<=result;
chainin_reg<=chainin; 
end
end

wire [4:0] flags1,flags2,flags3,flags4; 

FPMult_16_dspchain inst1(.clk(clk),.rst(reset),.a(top_a_reg),.b(top_b_reg),.flags(flags1),.result(r1)); 
FPMult_16_dspchain inst2(.clk(clk),.rst(reset),.a(bot_a_reg),.b(bot_b_reg),.flags(flags2),.result(r2));
FPAddSub_single_dspchain inst3(.clk(clk),.rst(reset),.a(r1),.b(r2),.flags(flags3),.operation(1'b1),.result(r3));
FPAddSub_single_dspchain inst4(.clk(clk),.rst(reset),.a(r3),.b(chainin),.flags(flags4),.operation(1'b1),.result(result));
assign chainout = result; 
endmodule
//`endif

//`timescale 1ns / 1ps


// IEEE Half Precision => 5 = 5, 10 = 10



//`define IEEE_COMPLIANCE 1


//////////////////////////////////////////////////////////////////////////////////
//
// Module Name:    FPMult
//
//////////////////////////////////////////////////////////////////////////////////

module FPMult_16_dspchain(
		clk,
		rst,
		a,
		b,
		result,
		flags
    );
	
	// Input Ports
	input clk ;							// Clock
	input rst ;							// Reset signal
	input [16-1:0] a;						// Input A, a 32-bit floating point number
	input [16-1:0] b;						// Input B, a 32-bit floating point number
	
	// Output ports
	output [32-1:0] result ;					// Product, result of the operation, 32-bit FP number
	output [4:0] flags ;						// Flags indicating exceptions according to IEEE754
	
	// Internal signals
	wire [32-1:0] Z_int ;					// Product, result of the operation, 32-bit FP number
	wire [4:0] Flags_int ;						// Flags indicating exceptions according to IEEE754
	
	wire Sa ;							// A's sign
	wire Sb ;							// B's sign
	wire Sp ;							// Product sign
	wire [5-1:0] Ea ;					// A's 5
	wire [5-1:0] Eb ;					// B's 5
	wire [2*10+1:0] Mp ;					// Product 10
	wire [4:0] InputExc ;						// Exceptions in inputs
	wire [23-1:0] NormM ;					// Normalized 10
	wire [8:0] NormE ;					// Normalized 5
	wire [23:0] RoundM ;					// Normalized 10
	wire [8:0] RoundE ;					// Normalized 5
	wire [23:0] RoundMP ;					// Normalized 10
	wire [8:0] RoundEP ;					// Normalized 5
	wire GRS ;

	//reg [63:0] pipe_0;						// Pipeline register Input->Prep
	reg [2*16-1:0] pipe_0;					// Pipeline register Input->Prep

	//reg [92:0] pipe_1;						// Pipeline register Prep->Execute
	//reg [3*10+2*5+7:0] pipe_1;			// Pipeline register Prep->Execute
	reg [3*10+2*5+18:0] pipe_1;

	//reg [38:0] pipe_2;						// Pipeline register Execute->Normalize
	reg [23+8+7:0] pipe_2;				// Pipeline register Execute->Normalize

	//reg [72:0] pipe_3;						// Pipeline register Normalize->Round
	reg [2*23+2*8+10:0] pipe_3;			// Pipeline register Normalize->Round

	//reg [36:0] pipe_4;						// Pipeline register Round->Output
	reg [32+4:0] pipe_4;					// Pipeline register Round->Output
	
	assign result = pipe_4[32+4:5] ;
	assign flags = pipe_4[4:0] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPMult_PrepModule_dspchain PrepModule(clk, rst, pipe_0[2*16-1:16], pipe_0[16-1:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10+1:0], InputExc[4:0]) ;

	// Perform (unsigned) 10 multiplication
	FPMult_ExecuteModule_dspchain ExecuteModule(pipe_1[3*10+5*2+7:2*10+2*5+8], pipe_1[2*10+2*5+7:2*10+7], pipe_1[2*10+6:5], pipe_1[2*10+2*5+6:2*10+5+7], pipe_1[2*10+5+6:2*10+7], pipe_1[2*10+2*5+8], pipe_1[2*10+2*5+7], Sp, NormE[8:0], NormM[23-1:0], GRS) ;

	// Round result and if necessary, perform a second (post-rounding) normalization step
	FPMult_NormalizeModule_dspchain NormalizeModule(pipe_2[23-1:0], pipe_2[23+8:23], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]) ;		

	// Round result and if necessary, perform a second (post-rounding) normalization step
	//FPMult_RoundModule RoundModule(pipe_3[47:24], pipe_3[23:0], pipe_3[65:57], pipe_3[56:48], pipe_3[66], pipe_3[67], pipe_3[72:68], Z_int[31:0], Flags_int[4:0]) ;		
	FPMult_RoundModule_dspchain RoundModule(pipe_3[2*23+1:23+1], pipe_3[23:0], pipe_3[2*8+2*23+3:2*23+8+3], pipe_3[2*23+8+2:2*23+2], pipe_3[2*23+2*8+4], pipe_3[2*23+2*8+5], pipe_3[2*23+2*8+10:2*23+2*8+6], Z_int[32-1:0], Flags_int[4:0]) ;		


//adding always@ (*) instead of posedge clock to make design combinational
	always @ (*) begin	
		if(rst) begin
			pipe_0 = 0;
			pipe_1 = 0;
			pipe_2 = 0; 
			pipe_3 = 0;
			pipe_4 = 0;
		end 
		else begin		
			/* PIPE 0
				[2*16-1:16] A
				[16-1:0] B
			*/
                       pipe_0 = {a, b} ;


			/* PIPE 1
				[2*5+3*10 + 18: 2*5+2*10 + 18] //pipe_0[16+10-1:16] , 10 of A
				[2*5+2*10 + 17 :2*5+2*10 + 9] // pipe_0[8:0]
				[2*5+2*10 + 8] Sa
				[2*5+2*10 + 7] Sb
				[2*5+2*10 + 6:5+2*10+7] Ea
				[5 +2*10+6:2*10+7] Eb
				[2*10+1+5:5] Mp
				[4:0] InputExc
			*/
			//pipe_1 <= {pipe_0[16+10-1:16], pipe_0[10_MUL_SPLIT_LSB-1:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10-1:0], InputExc[4:0]} ;
			pipe_1 = {pipe_0[16+10-1:16], pipe_0[8:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10+1:0], InputExc[4:0]} ;
			
			/* PIPE 2
				[8 + 23 + 7:8 + 23 + 3] InputExc
				[8 + 23 + 2] GRS
				[8 + 23 + 1] Sp
				[8 + 23:23] NormE
				[23-1:0] NormM
			*/
			pipe_2 = {pipe_1[4:0], GRS, Sp, NormE[8:0], NormM[23-1:0]} ;
			/* PIPE 3
				[2*8+2*23+10:2*8+2*23+6] InputExc
				[2*8+2*23+5] GRS
				[2*8+2*23+4] Sp	
				[2*8+2*23+3:8+2*23+3] RoundE
				[8+2*23+2:2*23+2] RoundEP
				[2*23+1:23+1] RoundM
				[23:0] RoundMP
			*/
			pipe_3 = {pipe_2[8 + 23 + 7:8 + 23 + 1], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]} ;
			/* PIPE 4
				[16+4:5] Z
				[4:0] Flags
			*/				
			pipe_4 = {Z_int[32-1:0], Flags_int[4:0]} ;
		end
	end
		
endmodule



module FPMult_PrepModule_dspchain (
		clk,
		rst,
		a,
		b,
		Sa,
		Sb,
		Ea,
		Eb,
		Mp,
		InputExc
	);
	
	// Input ports
	input clk ;
	input rst ;
	input [16-1:0] a ;								// Input A, a 32-bit floating point number
	input [16-1:0] b ;								// Input B, a 32-bit floating point number
	
	// Output ports
	output Sa ;										// A's sign
	output Sb ;										// B's sign
	output [5-1:0] Ea ;								// A's 5
	output [5-1:0] Eb ;								// B's 5
	output [2*10+1:0] Mp ;							// 10 product
	output [4:0] InputExc ;						// Input numbers are exceptions
	
	// Internal signals							// If signal is high...
	wire ANaN ;										// A is a signalling NaN
	wire BNaN ;										// B is a signalling NaN
	wire AInf ;										// A is infinity
	wire BInf ;										// B is infinity
    wire [10-1:0] Ma;
    wire [10-1:0] Mb;
	
	assign ANaN = &(a[16-2:10]) &  |(a[16-2:10]) ;			// All one 5 and not all zero 10 - NaN
	assign BNaN = &(b[16-2:10]) &  |(b[10-1:0]);			// All one 5 and not all zero 10 - NaN
	assign AInf = &(a[16-2:10]) & ~|(a[16-2:10]) ;		// All one 5 and all zero 10 - Infinity
	assign BInf = &(b[16-2:10]) & ~|(b[16-2:10]) ;		// All one 5 and all zero 10 - Infinity
	
	// Check for any exceptions and put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	//assign InputExc = {(ANaN | ANaN | BNaN |BNaN), ANaN, ANaN, BNaN,BNaN} ;
	
	// Take input numbers apart
	assign Sa = a[16-1] ;							// A's sign
	assign Sb = b[16-1] ;							// B's sign
	assign Ea = a[16-2:10];						// Store A's 5 in Ea, unless A is an exception
	assign Eb = b[16-2:10];						// Store B's 5 in Eb, unless B is an exception	
//    assign Ma = a[10_MSB:10_LSB];
  //  assign Mb = b[10_MSB:10_LSB];
	

	// Actual 10 multiplication occurs here
	//assign Mp = ({4'b0001, a[10-1:0]}*{4'b0001, b[10-1:9]}) ;
	assign Mp = ({1'b1,a[10-1:0]}*{1'b1, b[10-1:0]}) ;

	
    //We multiply part of the 10 here
    //Full 10 of A
    //Bits 10_MUL_SPLIT_MSB:10_MUL_SPLIT_LSB of B
   // wire [`ACTUAL_10-1:0] inp_A;
   // wire [`ACTUAL_10-1:0] inp_B;
   // assign inp_A = {1'b1, Ma};
   // assign inp_B = {{(10-(10_MUL_SPLIT_MSB-10_MUL_SPLIT_LSB+1)){1'b0}}, 1'b1, Mb[10_MUL_SPLIT_MSB:10_MUL_SPLIT_LSB]};
   // DW02_mult #(`ACTUAL_10,`ACTUAL_10) u_mult(.A(inp_A), .B(inp_B), .TC(1'b0), .PRODUCT(Mp));
endmodule


module FPMult_ExecuteModule_dspchain(
		a,
		b,
		MpC,
		Ea,
		Eb,
		Sa,
		Sb,
		Sp,
		NormE,
		NormM,
		GRS
    );

	// Input ports
	input [10-1:0] a ;
	input [2*5:0] b ;
	input [2*10+1:0] MpC ;
	input [5-1:0] Ea ;						// A's 5
	input [5-1:0] Eb ;						// B's 5
	input Sa ;								// A's sign
	input Sb ;								// B's sign
	
	// Output ports
	output Sp ;								// Product sign
	output [8:0] NormE ;													// Normalized 5
	output [23-1:0] NormM ;												// Normalized 10
	output GRS ;
	
	wire [2*10+1:0] Mp ;
	
	assign Sp = (Sa ^ Sb) ;												// Equal signs give a positive product
	
   // wire [`ACTUAL_10-1:0] inp_a;
   // wire [`ACTUAL_10-1:0] inp_b;
   // assign inp_a = {1'b1, a};
   // assign inp_b = {{(10-10_MUL_SPLIT_LSB){1'b0}}, 1'b0, b};
   // DW02_mult #(`ACTUAL_10,`ACTUAL_10) u_mult(.A(inp_a), .B(inp_b), .TC(1'b0), .PRODUCT(Mp_temp));
   // DW01_add #(2*`ACTUAL_10) u_add(.A(Mp_temp), .B(MpC<<10_MUL_SPLIT_LSB), .CI(1'b0), .SUM(Mp), .CO());

	//assign Mp = (MpC<<(2*5+1)) + ({4'b0001, a[10-1:0]}*{1'b0, b[2*5:0]}) ;
	assign Mp = MpC;


	assign NormM = (Mp[2*10+1] ? Mp[2*10:0] : Mp[2*10-1:0]); 	// Check for overflow
	assign NormE = (Ea + Eb + Mp[2*10+1]);								// If so, increment 5
	
	assign GRS = ((Mp[10]&(Mp[10+1]))|(|Mp[10-1:0])) ;
	
endmodule

module FPMult_NormalizeModule_dspchain(
		NormM,
		NormE,
		RoundE,
		RoundEP,
		RoundM,
		RoundMP
    );

	// Input Ports
	input [23-1:0] NormM ;									// Normalized 10
	input [8:0] NormE ;									// Normalized 5

	// Output Ports
	output [8:0] RoundE ;
	output [8:0] RoundEP ;
	output [23:0] RoundM ;
	output [23:0] RoundMP ; 
	
// 5 = 5 
// 5 -1 = 4
// NEED to subtract 2^4 -1 = 15

wire [8-1 : 0] bias;

assign bias =  ((1<< (8 -1)) -1);

	assign RoundE = NormE - 9'd15 - 9'd15 + 9'd127 ;
	assign RoundEP = NormE - 9'd15 - 9'd15 + 9'd127 ;
	assign RoundM = NormM ;
	assign RoundMP = NormM ;

endmodule

module FPMult_RoundModule_dspchain(
		RoundM,
		RoundMP,
		RoundE,
		RoundEP,
		Sp,
		GRS,
		InputExc,
		Z,
		Flags
    );

	// Input Ports
	input [23:0] RoundM ;									// Normalized 10
	input [23:0] RoundMP ;									// Normalized 5
	input [8:0] RoundE ;									// Normalized 10 + 1
	input [8:0] RoundEP ;									// Normalized 5 + 1
	input Sp ;												// Product sign
	input GRS ;
	input [4:0] InputExc ;
	
	// Output Ports
	output [32-1:0] Z ;										// Final product
	output [4:0] Flags ;
	
	// Internal Signals
	wire [8:0] FinalE ;									// Rounded 5
	wire [23:0] FinalM;
	wire [23:0] PreShiftM;
	
	assign PreShiftM = GRS ? RoundMP : RoundM ;	// Round up if R and (G or S)
	
	// Post rounding normalization (potential one bit shift> use shifted 10 if there is overflow)
	assign FinalM = (PreShiftM[23] ? {1'b0, PreShiftM[23:1]} : PreShiftM[23:0]) ;
	assign FinalE = (PreShiftM[23] ? RoundEP : RoundE) ; // Increment 5 if a shift was done
	
	
	assign Z = {Sp, FinalE[8-1:0], FinalM[21-1:0], 2'b0} ;   // Putting the pieces together
	assign Flags = InputExc[4:0];

endmodule


module FPAddSub_single_dspchain(
		clk,
		rst,
		a,
		b,
		operation,
		result,
		flags
	);

// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [31:0] a ;								// Input A, a 32-bit floating point number
	input [31:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [31:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754

	reg [68:0]pipe_1;
	reg [54:0]pipe_2;
	reg [45:0]pipe_3;


//internal module wires

//output ports
	wire Opout;
	wire Sa;
	wire Sb;
	wire MaxAB;
	wire [7:0] CExp;
	wire [4:0] Shift;
	wire [22:0] Mmax;
	wire [4:0] InputExc;
	wire [23:0] Mmin_3;

	wire [32:0] SumS_5 ;
	wire [4:0] Shift_1;							
	wire PSgn ;							
	wire Opr ;	
	
	wire [22:0] NormM ;				// Normalized mantissa
	wire [8:0] NormE ;					// Adjusted exponent
	wire ZeroSum ;						// Zero flag
	wire NegE ;							// Flag indicating negative exponent
	wire R ;								// Round bit
	wire S ;								// Final sticky bit
	wire FG ;

FPAddSub_a_dspchain M1(a,b,operation,Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3);

FpAddSub_b_dspchain M2(pipe_1[51:29],pipe_1[23:0],pipe_1[67],pipe_1[66],pipe_1[65],pipe_1[68],SumS_5,Shift_1,PSgn,Opr);

FPAddSub_c_dspchain M3(pipe_2[54:22],pipe_2[21:17],pipe_2[16:9],NormM,NormE,ZeroSum,NegE,R,S,FG);

FPAddSub_d_dspchain M4(pipe_3[13],pipe_3[22:14],pipe_3[45:23],pipe_3[11],pipe_3[10],pipe_3[9],pipe_3[8],pipe_3[7],pipe_3[6],pipe_3[5],pipe_3[12],pipe_3[4:0],result,flags );


always @ (posedge clk) begin	
		if(rst) begin
			pipe_1 <= 0;
			pipe_2 <= 0;
			pipe_3 <= 0;
		end 
		else begin
/*
pipe_1:
	[68] Opout;
	[67] Sa;
	[66] Sb;
	[65] MaxAB;
	[64:57] CExp;
	[56:52] Shift;
	[51:29] Mmax;
	[28:24] InputExc;
	[23:0] Mmin_3;	
*/

pipe_1 <= {Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3};

/*
pipe_2:
	[54:22]SumS_5;
	[21:17]Shift;
	[16:9]CExp;	
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_2 <= {SumS_5,Shift_1,pipe_1[64:57], pipe_1[67], pipe_1[66], pipe_1[68], pipe_1[65], pipe_1[28:24] };

/*
pipe_3:
	[45:23] NormM ;				
	[22:14] NormE ;					
	[13]ZeroSum ;						
	[12]NegE ;							
	[11]R ;								
	[10]S ;								
	[9]FG ;
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_3 <= {NormM,NormE,ZeroSum,NegE,R,S,FG, pipe_2[8], pipe_2[7], pipe_2[6], pipe_2[5], pipe_2[4:0] };

end
end

endmodule

// Prealign + Align + Shift 1 + Shift 2
module FPAddSub_a_dspchain(
		A,
		B,
		operation,
		Opout,
		Sa,
		Sb,
		MaxAB,
		CExp,
		Shift,
		Mmax,
		InputExc,
		Mmin_3
		
		
	);
	
	// Input ports
	input [31:0] A ;										// Input A, a 32-bit floating point number
	input [31:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	//output ports
	output Opout;
	output Sa;
	output Sb;
	output MaxAB;
	output [7:0] CExp;
	output [4:0] Shift;
	output [22:0] Mmax;
	output [4:0] InputExc;
	output [23:0] Mmin_3;	
							
	wire [9:0] ShiftDet ;							
	wire [30:0] Aout ;
	wire [30:0] Bout ;
	

	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [7:0] DAB ;										// ExpA - ExpB					
	wire [7:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[30:23]) & |(A[22:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[30:23]) & |(B[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[30:23]) & ~|(A[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[30:23]) & ~|(B[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
  assign DAB = (A[30:23] + ~(B[30:23]) + 1) ;
	assign DBA = (B[30:23] + ~(A[30:23]) + 1) ;

	assign Sa = A[31] ;									// A's sign bit
	assign Sb = B[31] ;									// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[30:0] ;
	assign Bout = B[30:0] ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Output ports
													// Number of steps to smaller mantissa shift right
	wire [22:0] Mmin_1 ;							// Smaller mantissa 
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (Aout[30:0] < Bout[30:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[9:5] : ShiftDet[4:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin_1 = MaxAB ? Aout[22:0] : Bout[22:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? Bout[22:0]: Aout[22:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? Bout[30:23] : Aout[30:23]) ;	

// Input ports
					// Smaller mantissa after 16|12|8|4 shift
	wire [2:0] Shift_1 ;						// Shift amount
	
	assign Shift_1 = Shift [4:2];

	wire [23:0] Mmin_2 ;						// The smaller mantissa
	
	// Internal signals
	reg	  [23:0]		Lvl1;
	reg	  [23:0]		Lvl2;
	wire    [47:0]    Stage1;	
	integer           i;                // Loop variable
	
	always @(*) begin						
		// Rotate by 16?
		Lvl1 <= Shift_1[2] ? {17'b00000000000000001, Mmin_1[22:16]} : {1'b1, Mmin_1}; 
	end
	
	assign Stage1 = {Lvl1, Lvl1};
	
	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift_1[1:0])
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[23:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[23:19] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[23:15] <= 0; end
			// Rotate by 12	
			2'b11:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[23:11] <= 0; end
	  endcase
	end
	
	// Assign output to next shift stage
	assign Mmin_2 = Lvl2;
								// Smaller mantissa after 16|12|8|4 shift
	wire [1:0] Shift_2 ;						// Shift amount
	
	assign Shift_2 =Shift  [1:0] ;
					// The smaller mantissa
	
	// Internal Signal
	reg	  [23:0]		Lvl3;
	wire    [47:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {Mmin_2, Mmin_2};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_2[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[23:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[23] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[23:22] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[23:21] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin_3 = Lvl3;	

	
endmodule

module FpAddSub_b_dspchain(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		SumS_5,
		Shift,
		PSgn,
		Opr
);
	input [22:0] Mmax ;					// The larger mantissa
	input [23:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	wire [32:0] Sum ;	
						// Output ports
	output [32:0] SumS_5 ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount				// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation

	// Perform effective operation
	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, 8'b00000000} - {Mmin, 8'b00000000}) : ({1'b1, Mmax, 8'b00000000} + {Mmin, 8'b00000000}) ;
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

		// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[32] ? 5'b00000 :	 
		Sum[31] ? 5'b00001 : 
		Sum[30] ? 5'b00010 : 
		Sum[29] ? 5'b00011 : 
		Sum[28] ? 5'b00100 : 
		Sum[27] ? 5'b00101 : 
		Sum[26] ? 5'b00110 : 
		Sum[25] ? 5'b00111 :
		Sum[24] ? 5'b01000 :
		Sum[23] ? 5'b01001 :
		Sum[22] ? 5'b01010 :
		Sum[21] ? 5'b01011 :
		Sum[20] ? 5'b01100 :
		Sum[19] ? 5'b01101 :
		Sum[18] ? 5'b01110 :
		Sum[17] ? 5'b01111 :
		Sum[16] ? 5'b10000 :
		Sum[15] ? 5'b10001 :
		Sum[14] ? 5'b10010 :
		Sum[13] ? 5'b10011 :
		Sum[12] ? 5'b10100 :
		Sum[11] ? 5'b10101 :
		Sum[10] ? 5'b10110 :
		Sum[9] ? 5'b10111 :
		Sum[8] ? 5'b11000 :
		Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [32:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[16:0], 16'b0000000000000000} : Sum; 
	end
	
	// Assign outputs
	assign SumS_5 = Lvl1;	

endmodule

module FPAddSub_c_dspchain(
		SumS_5,
		Shift,
		CExp,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [32:0] SumS_5 ;						// Smaller mantissa after 16|12|8|4 shift
	
	input [4:0] Shift ;						// Shift amount
	
// Input ports
	
	input [7:0] CExp ;
	

	// Output ports
	output [22:0] NormM ;				// Normalized mantissa
	output [8:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;


	wire [3:0]Shift_1;
	assign Shift_1 = Shift [3:0];
	// Output ports
	wire [32:0] SumS_7 ;						// The smaller mantissa
	
	reg	  [32:0]		Lvl2;
	wire    [65:0]    Stage1;	
	reg	  [32:0]		Lvl3;
	wire    [65:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {SumS_5, SumS_5};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[32:0];       		
			// Rotate by 4
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_1[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[32:0];
			// Rotate by 1
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign SumS_7 = Lvl3;						// Take out smaller mantissa



	
	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [8:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [8:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = SumS_7[32] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|SumS_7 ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[8] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = SumS_7[31:9] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = SumS_7[8] ; 
	assign R = SumS_7[7] ;
	assign S = |SumS_7[6:0] ;		
	
endmodule

module FPAddSub_d_dspchain(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		NegE,
		InputExc,
		P,
		Flags 
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [8:0] NormE ;				// Normalized exponent
	input [22:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	

	input NegE ;						// Negative exponent?
	input [4:0] InputExc ;					// Exceptions in inputs A and B

	// Output ports
	output [31:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// 
	wire [31:0] Z ;					// Final result
	wire EOF ;
	
	// Internal signals
	wire [23:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [22:0] RoundM ;				// The final rounded sum
	wire [8:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	wire FSgn;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[22:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[23] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? 8'b00000000 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[7:0], RoundM[22:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[8];

/////////////////////////////////////////////////////////////////////////////////////////////////////////



	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[30:23]) & ~|(Z[30:23]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule

`endif 


module fifo_512_60bit
	#(parameter dw=60,
	  parameter aw=9)
	(clk, rst, clr, din, we, dout, re,
	full, empty);

parameter max_size = 1<<aw;

input 			clk, rst, clr;
input 	[dw-1:0]	din;
input 			we;
output	[dw-1:0]	dout;
input 	wire		re;
output			full;
output			empty;

////////////////////////////////////////////////////////////////////
//
// Local Wires
//
wire 	[dw-1:0]	din_nc;
wire 	[dw-1:0]	out_nc;
reg		[aw-1:0]	wp;
wire	[aw-1:0]	wp_pl1;
reg		[aw-1:0]	rp;
wire	[aw-1:0]	rp_pl1;
reg					gb;

////////////////////////////////////////////////////////////////////
//
// Memory Block
//
dpram_512_60bit #(
	.AWIDTH(aw),
	.DWIDTH(dw)
	) u0 (
	.clk(clk),
	.address_a(rp),
	.wren_a(0),
	.data_a(din_nc),
	.out_a(dout),
	.address_b(wp),
	.wren_b(we),
	.data_b(din),
	.out_b(out_nc)
);


////////////////////////////////////////////////////////////////////
//
// Misc Logic
//

always @(posedge clk or posedge rst)
	if(rst)	wp <= {aw{1'b0}};
	else
	if(clr)		wp <= {aw{1'b0}};
	else
	if(we)		wp <= wp_pl1;

assign wp_pl1 = wp + { {aw-1{1'b0}}, 1'b1};

always @(posedge clk or posedge rst)
	if(rst)		rp <= {aw{1'b0}};
	else
	if(clr)		rp <= {aw{1'b0}};
	else
	if(re)		rp <= rp_pl1;

assign rp_pl1 = rp + { {aw-1{1'b0}}, 1'b1};

////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//

assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);

// Guard Bit ...
always @(posedge clk or posedge rst)
	if(rst)						gb <= 1'b0;
	else
	if(clr)						gb <= 1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <= 1'b1;
	else
	if(re)						gb <= 1'b0;

endmodule

module dpram_512_60bit #(
	parameter DWIDTH = 60,
	parameter AWIDTH = 9
  )
  (
	clk,
	address_a,
	address_b,
	wren_a,
	wren_b,
	data_a,
	data_b,
	out_a,
	out_b
);

parameter NUM_WORDS=1<<AWIDTH;

input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

	reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];

	always @ (posedge clk) begin
		if (wren_a) begin
			ram[address_a] <= data_a;
		end
		else begin
			out_a <= ram[address_a];
		end
	end
	  
	always @ (posedge clk) begin 
		if (wren_b) begin
			ram[address_b] <= data_b;
		end 
		else begin
			out_b <= ram[address_b];
		end
	end

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

	dual_port_ram u_dual_port_ram(
	.addr1(address_a),
	.we1(wren_a),
	.data1(data_a),
	.out1(out_a),
	.addr2(address_b),
	.we2(wren_b),
	.data2(data_b),
	.out2(out_b),
	.clk(clk)
	);

`endif

endmodule

module fifo_256_40bit
	#(parameter dw=40,
	  parameter aw=8)
	(clk, rst, clr, din, we, dout, re,
	full, empty);

parameter max_size = 1<<aw;

input 			clk, rst, clr;
input 	[dw-1:0]	din;
input 			we;
output	[dw-1:0]	dout;
input 	wire		re;
output			full;
output			empty;

////////////////////////////////////////////////////////////////////
//
// Local Wires
//
wire 	[dw-1:0]	din_nc;
wire 	[dw-1:0]	out_nc;
reg		[aw-1:0]	wp;
wire	[aw-1:0]	wp_pl1;
reg		[aw-1:0]	rp;
wire	[aw-1:0]	rp_pl1;
reg					gb;

////////////////////////////////////////////////////////////////////
//
// Memory Block
//
dpram_256_40bit #(
	.AWIDTH(aw),
	.DWIDTH(dw)
	) u0 (
	.clk(clk),
	.address_a(rp),
	.wren_a(0),
	.data_a(din_nc),
	.out_a(dout),
	.address_b(wp),
	.wren_b(we),
	.data_b(din),
	.out_b(out_nc)
);


////////////////////////////////////////////////////////////////////
//
// Misc Logic
//

always @(posedge clk or posedge rst)
	if(rst)	wp <= {aw{1'b0}};
	else
	if(clr)		wp <= {aw{1'b0}};
	else
	if(we)		wp <= wp_pl1;

assign wp_pl1 = wp + { {aw-1{1'b0}}, 1'b1};

always @(posedge clk or posedge rst)
	if(rst)		rp <= {aw{1'b0}};
	else
	if(clr)		rp <= {aw{1'b0}};
	else
	if(re)		rp <= rp_pl1;

assign rp_pl1 = rp + { {aw-1{1'b0}}, 1'b1};

////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//

assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);

// Guard Bit ...
always @(posedge clk or posedge rst)
	if(rst)						gb <= 1'b0;
	else
	if(clr)						gb <= 1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <= 1'b1;
	else
	if(re)						gb <= 1'b0;

endmodule

module dpram_256_40bit #(
	parameter DWIDTH = 40,
	parameter AWIDTH = 8
  )
  (
	clk,
	address_a,
	address_b,
	wren_a,
	wren_b,
	data_a,
	data_b,
	out_a,
	out_b
);

parameter NUM_WORDS=1<<AWIDTH;

input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

	reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];

	always @ (posedge clk) begin
		if (wren_a) begin
			ram[address_a] <= data_a;
		end
		else begin
			out_a <= ram[address_a];
		end
	end
	  
	always @ (posedge clk) begin 
		if (wren_b) begin
			ram[address_b] <= data_b;
		end 
		else begin
			out_b <= ram[address_b];
		end
	end

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;


	dual_port_ram u_dual_port_ram(
	.addr1(address_a),
	.we1(wren_a),
	.data1(data_a),
	.out1(out_a),
	.addr2(address_b),
	.we2(wren_b),
	.data2(data_b),
	.out2(out_b),
	.clk(clk)
	);

`endif

endmodule
module tensor_block(
	clk,
	reset,
	
	data_in,
	cascade_in,
	acc0_in,
	acc1_in,
	acc2_in,
	accumulator_input1_select,

	out0,
	out1,
	out2,
	cascade_out,
	acc0_out,
	acc1_out,
	acc2_out,

	mux1_select,
	dot_unit_input_1_enable,
	bank0_data_in_enable,
	bank1_data_in_enable,
	cascade_out_select,
	dot_unit_input_2_select

	);

input 	[79:0] data_in;
input	[79:0] cascade_in;
input	[31:0] acc0_in;
input	[31:0] acc1_in;
input	[31:0] acc2_in;
input 	[2:0] accumulator_input1_select;


output	[24:0] out0;
output	[24:0] out1;
output	[24:0] out2;
output	[79:0] cascade_out;
output	[31:0] acc0_out;
output	[31:0] acc1_out;
output	[31:0] acc2_out;

//Inputs to take into account
input clk;
input reset;

// Logic to be created for 
input mux1_select;
input dot_unit_input_1_enable;
input bank0_data_in_enable;
input bank1_data_in_enable;
input cascade_out_select;
input dot_unit_input_2_select;


wire [79:0]mux1_out;
assign mux1_out = mux1_select ? cascade_in : data_in;

reg [79:0]dot_unit_input_1;

// D Flip Flop with reset and enable
always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) dot_unit_input_1 <= 0;
	else if (dot_unit_input_1_enable) dot_unit_input_1 <= data_in;
end

// Register Bank 0 
reg[79:0] bank0_reg0;
reg[79:0] bank0_reg1;
reg[79:0] bank0_reg2;

always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) begin
		bank0_reg0 <= 0;
		bank0_reg1 <= 0;
		bank0_reg2 <= 0;
	end
	else if (bank0_data_in_enable) begin
		bank0_reg0 <= mux1_out;
		bank0_reg1 <= bank0_reg0;
		bank0_reg2 <= bank0_reg1;
	end
end

// Register Bank 1 
reg[79:0] bank1_reg0;
reg[79:0] bank1_reg1;
reg[79:0] bank1_reg2;

always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) begin
		bank1_reg0 <= 0;
		bank1_reg1 <= 0;
		bank1_reg2 <= 0;
	end
	else if (bank1_data_in_enable) begin
		bank1_reg0 <= mux1_out;
		bank1_reg1 <= bank0_reg0;
		bank1_reg2 <= bank0_reg1;
	end
end

// Output cascade out
assign cascade_out = cascade_out_select ? bank1_reg2 : bank0_reg2;

// Providing second input to all 3 dot product units
wire [79:0]dot_unit_input_2_0;
wire [79:0]dot_unit_input_2_1;
wire [79:0]dot_unit_input_2_2;

assign dot_unit_input_2_0 = dot_unit_input_2_select ? bank1_reg0 : bank0_reg0;
assign dot_unit_input_2_1 = dot_unit_input_2_select ? bank1_reg1 : bank0_reg1;
assign dot_unit_input_2_2 = dot_unit_input_2_select ? bank1_reg2 : bank0_reg2;

wire [19:0] dot_unit_output_0;
wire [19:0] dot_unit_output_1;
wire [19:0] dot_unit_output_2;

dot_product_unit dot_unit0 (dot_unit_input_1, dot_unit_input_2_0, dot_unit_output_0,clk);
dot_product_unit dot_unit1 (dot_unit_input_1, dot_unit_input_2_1, dot_unit_output_1,clk);
dot_product_unit dot_unit2 (dot_unit_input_1, dot_unit_input_2_2, dot_unit_output_2,clk);

// Flopping after dot product compute
reg [19:0] dot_unit_output_0_flopped;
reg [19:0] dot_unit_output_1_flopped;
reg [19:0] dot_unit_output_2_flopped;

always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) begin
		dot_unit_output_0_flopped <= 0;
		dot_unit_output_1_flopped <= 0;
		dot_unit_output_2_flopped <= 0;
	end
	else begin
		dot_unit_output_0_flopped <= dot_unit_output_0;
		dot_unit_output_1_flopped <= dot_unit_output_1;
		dot_unit_output_2_flopped <= dot_unit_output_2;
	end
end

wire [31:0] accumulator_unit0_input1;
wire [31:0] accumulator_unit1_input1;
wire [31:0] accumulator_unit2_input1;

wire [31:0] accumulator_unit_output_0;
wire [31:0] accumulator_unit_output_1;
wire [31:0] accumulator_unit_output_2;

reg [31:0] accumulator_unit_output_0_flopped;
reg [31:0] accumulator_unit_output_1_flopped;
reg [31:0] accumulator_unit_output_2_flopped;

reg [31:0] acc0_in_flopped;
reg [31:0] acc1_in_flopped;
reg [31:0] acc2_in_flopped;

// 3 mux's for selecting acc_in or acc_out_flopped
assign accumulator_unit0_input1 = accumulator_input1_select[0] ?  accumulator_unit_output_0_flopped : acc0_in_flopped;
assign accumulator_unit1_input1 = accumulator_input1_select[1] ?  accumulator_unit_output_1_flopped : acc1_in_flopped;
assign accumulator_unit2_input1 = accumulator_input1_select[2] ?  accumulator_unit_output_2_flopped : acc2_in_flopped;

// Flopping the accumulator outputs and acc_in 
always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) begin
		accumulator_unit_output_0_flopped <= 0;
		accumulator_unit_output_1_flopped <= 0;
		accumulator_unit_output_2_flopped <= 0;
		acc0_in_flopped <= 0;
		acc1_in_flopped <= 0;
		acc2_in_flopped <= 0;
	end
	else begin
		accumulator_unit_output_0_flopped <= accumulator_unit_output_0;
		accumulator_unit_output_1_flopped <= accumulator_unit_output_1;
		accumulator_unit_output_2_flopped <= accumulator_unit_output_2;
		acc0_in_flopped <= acc0_in;
		acc1_in_flopped <= acc1_in;
		acc2_in_flopped <= acc2_in;
	end
end

// Accumulator units
accumulator acc_unit0 (dot_unit_output_0_flopped, accumulator_unit0_input1, accumulator_unit_output_0 );
accumulator acc_unit1 (dot_unit_output_1_flopped, accumulator_unit1_input1, accumulator_unit_output_1 );
accumulator acc_unit2 (dot_unit_output_2_flopped, accumulator_unit2_input1, accumulator_unit_output_2 );

assign acc0_out = accumulator_unit_output_0;
assign acc1_out = accumulator_unit_output_1;
assign acc2_out = accumulator_unit_output_2;

//Taking the top 25 bits from the 32 bit accumulation number
assign out0= accumulator_unit_output_0[31:7];
assign out1= accumulator_unit_output_1[31:7];
assign out2= accumulator_unit_output_2[31:7];

endmodule

module dot_product_unit (
	data_in_1,
	data_in_2,
	data_out,
  clk
	);

input clk;
input [79:0] data_in_1;
input [79:0] data_in_2;
output reg [19:0] data_out;

wire [7:0] mult1_in1;
wire [7:0] mult1_in2;
reg [15:0] mult1_out;
wire [7:0] mult2_in1;
wire [7:0] mult2_in2;
reg [15:0] mult2_out;
wire [7:0] mult3_in1;
wire [7:0] mult3_in2;
reg [15:0] mult3_out;
wire [7:0] mult4_in1;
wire [7:0] mult4_in2;
reg [15:0] mult4_out;
wire [7:0] mult5_in1;
wire [7:0] mult5_in2;
reg [15:0] mult5_out;
wire [7:0] mult6_in1;
wire [7:0] mult6_in2;
reg [15:0] mult6_out;
wire [7:0] mult7_in1;
wire [7:0] mult7_in2;
reg [15:0] mult7_out;
wire [7:0] mult8_in1;
wire [7:0] mult8_in2;
reg [15:0] mult8_out;
wire [7:0] mult9_in1;
wire [7:0] mult9_in2;
reg [15:0] mult9_out;
wire [7:0] mult10_in1;
wire [7:0] mult10_in2;
reg [15:0] mult10_out;

assign mult1_in1 = data_in_1[7:0];
assign mult1_in2 = data_in_2[7:0];

assign mult2_in1 = data_in_1[15:8];
assign mult2_in2 = data_in_2[15:8];


assign mult3_in1 = data_in_1[23:16];
assign mult3_in2 = data_in_2[23:16];

assign mult4_in1 = data_in_1[31:24];
assign mult4_in2 = data_in_2[31:24];

assign mult5_in1 = data_in_1[39:32];
assign mult5_in2 = data_in_2[39:32];

assign mult6_in1 = data_in_1[47:40];
assign mult6_in2 = data_in_2[47:40];

assign mult7_in1 = data_in_1[55:48];
assign mult7_in2 = data_in_2[55:48];

assign mult8_in1 = data_in_1[63:56];
assign mult8_in2 = data_in_2[63:56];

assign mult9_in1 = data_in_1[71:64];
assign mult9_in2 = data_in_2[71:64];


assign mult10_in1 = data_in_1[79:72];
assign mult10_in2 = data_in_2[79:72];

always@(posedge clk) begin 
mult1_out <= mult1_in1 * mult1_in2;
mult2_out <= mult2_in1 * mult2_in2;
mult3_out <= mult3_in1 * mult3_in2;
mult4_out <= mult4_in1 * mult4_in2;
mult5_out <= mult5_in1 * mult5_in2;
mult6_out <= mult6_in1 * mult6_in2;
mult7_out <= mult7_in1 * mult7_in2;
mult8_out <= mult8_in1 * mult8_in2;
mult9_out <= mult9_in1 * mult9_in2;
mult10_out <= mult10_in1 * mult10_in2;
end



reg [16:0] s01,s02,s03,s04,s05;

always@(posedge clk) begin 
  s01<= mult1_out + mult2_out;
  s02<= mult3_out + mult4_out;
  s03<= mult5_out + mult6_out;
  s04<= mult7_out + mult8_out;
  s05<= mult9_out + mult10_out;
end

reg [17:0] s11,s12;

always@(posedge clk) begin 
s11<= s01 + s02;
s12<= s03 + s04; 
end

reg [18:0] s21;

always@(posedge clk) begin 
s21<= s11 + s12;
data_out <= s21 + s05; 
end



endmodule


module accumulator (
	input_accumlator_1,
	input_accumlator_2,
	output_accumlator
	);

input [19:0] input_accumlator_1;
input [31:0] input_accumlator_2;
output [31:0] output_accumlator;

assign output_accumlator = input_accumlator_1 + input_accumlator_2;

endmodule

module dsp_chain_4_int_sop_2 (clk,reset,ax1,ay1,bx1,by1,ax2,ay2,bx2,by2,ax3,ay3,bx3,by3,ax4,ay4,bx4,by4,result);

input clk; 
input reset; 
input [17:0] ax1, bx1, ax2, bx2, ax3, bx3, ax4, bx4; 
input [18:0] ay1, by1, ay2, by2, ay3, by3, ay4, by4; 
output reg [36:0] result; 

wire [36:0] chainout0, chainout1, chainout2, chainout3; 
wire [36:0] chainin0, chainin1, chainin2, chainin3; 
wire [36:0] resulta1, resulta2, resulta3, resulta4;

assign chainin0 = 37'd0;

int_sop_2_dspchain inst1 (.clk(clk),.reset(reset),.ax(ax1),.bx(bx1),.ay(ay1),.by(by1),.mode_sigs(11'd0),.chainin(chainin0),.resulta(resulta1),.chainout(chainout0));
int_sop_2_dspchain inst2 (.clk(clk),.reset(reset),.ax(ax2),.bx(bx2),.ay(ay2),.by(by2),.mode_sigs(11'd0),.chainin(chainout0),.resulta(resulta2),.chainout(chainout1));
int_sop_2_dspchain inst3 (.clk(clk),.reset(reset),.ax(ax3),.bx(bx3),.ay(ay3),.by(by3),.mode_sigs(11'd0),.chainin(chainout1),.resulta(resulta3),.chainout(chainout2));
int_sop_2_dspchain inst4 (.clk(clk),.reset(reset),.ax(ax4),.bx(bx4),.ay(ay4),.by(by4),.mode_sigs(11'd0),.chainin(chainout2),.resulta(resulta4),.chainout(chainout3));

assign result = resulta4;



endmodule 
module fifo_256_60bit
	#(parameter dw=60,
	  parameter aw=8)
	(clk, rst, clr, din, we, dout, re,
	full, empty);

parameter max_size = 1<<aw;

input 			clk, rst, clr;
input 	[dw-1:0]	din;
input 			we;
output	[dw-1:0]	dout;
input 	wire		re;
output			full;
output			empty;

////////////////////////////////////////////////////////////////////
//
// Local Wires
//
wire 	[dw-1:0]	din_nc;
wire 	[dw-1:0]	out_nc;
reg		[aw-1:0]	wp;
wire	[aw-1:0]	wp_pl1;
reg		[aw-1:0]	rp;
wire	[aw-1:0]	rp_pl1;
reg					gb;

////////////////////////////////////////////////////////////////////
//
// Memory Block
//
dpram_256_60bit #(
	.AWIDTH(aw),
	.DWIDTH(dw)
	) u0 (
	.clk(clk),
	.address_a(rp),
	.wren_a(0),
	.data_a(din_nc),
	.out_a(dout),
	.address_b(wp),
	.wren_b(we),
	.data_b(din),
	.out_b(out_nc)
);


////////////////////////////////////////////////////////////////////
//
// Misc Logic
//

always @(posedge clk or posedge rst)
	if(rst)	wp <= {aw{1'b0}};
	else
	if(clr)		wp <= {aw{1'b0}};
	else
	if(we)		wp <= wp_pl1;

assign wp_pl1 = wp + { {aw-1{1'b0}}, 1'b1};

always @(posedge clk or posedge rst)
	if(rst)		rp <= {aw{1'b0}};
	else
	if(clr)		rp <= {aw{1'b0}};
	else
	if(re)		rp <= rp_pl1;

assign rp_pl1 = rp + { {aw-1{1'b0}}, 1'b1};

////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//

assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);

// Guard Bit ...
always @(posedge clk or posedge rst)
	if(rst)						gb <= 1'b0;
	else
	if(clr)						gb <= 1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <= 1'b1;
	else
	if(re)						gb <= 1'b0;

endmodule

module dpram_256_60bit #(
	parameter DWIDTH = 60,
	parameter AWIDTH = 8
  )
  (
	clk,
	address_a,
	address_b,
	wren_a,
	wren_b,
	data_a,
	data_b,
	out_a,
	out_b
);

parameter NUM_WORDS=1<<AWIDTH;

input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

	reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];

	always @ (posedge clk) begin
		if (wren_a) begin
			ram[address_a] <= data_a;
		end
		else begin
			out_a <= ram[address_a];
		end
	end
	  
	always @ (posedge clk) begin 
		if (wren_b) begin
			ram[address_b] <= data_b;
		end 
		else begin
			out_b <= ram[address_b];
		end
	end

`else
defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

	dual_port_ram u_dual_port_ram(
	.addr1(address_a),
	.we1(wren_a),
	.data1(data_a),
	.out1(out_a),
	.addr2(address_b),
	.we2(wren_b),
	.data2(data_b),
	.out2(out_b),
	.clk(clk)
	);

`endif

endmodule

module fifo_512_40bit
	#(parameter dw=40,
	  parameter aw=9)
	(clk, rst, clr, din, we, dout, re,
	full, empty);

parameter max_size = 1<<aw;

input 			clk, rst, clr;
input 	[dw-1:0]	din;
input 			we;
output	[dw-1:0]	dout;
input 	wire		re;
output			full;
output			empty;

////////////////////////////////////////////////////////////////////
//
// Local Wires
//
wire 	[dw-1:0]	din_nc;
wire 	[dw-1:0]	out_nc;
reg		[aw-1:0]	wp;
wire	[aw-1:0]	wp_pl1;
reg		[aw-1:0]	rp;
wire	[aw-1:0]	rp_pl1;
reg					gb;

////////////////////////////////////////////////////////////////////
//
// Memory Block
//
dpram_512_40bit #(
	.AWIDTH(aw),
	.DWIDTH(dw)
	) u0 (
	.clk(clk),
	.address_a(rp),
	.wren_a(0),
	.data_a(din_nc),
	.out_a(dout),
	.address_b(wp),
	.wren_b(we),
	.data_b(din),
	.out_b(out_nc)
);


////////////////////////////////////////////////////////////////////
//
// Misc Logic
//

always @(posedge clk or posedge rst)
	if(rst)	wp <= {aw{1'b0}};
	else
	if(clr)		wp <= {aw{1'b0}};
	else
	if(we)		wp <= wp_pl1;

assign wp_pl1 = wp + { {aw-1{1'b0}}, 1'b1};

always @(posedge clk or posedge rst)
	if(rst)		rp <= {aw{1'b0}};
	else
	if(clr)		rp <= {aw{1'b0}};
	else
	if(re)		rp <= rp_pl1;

assign rp_pl1 = rp + { {aw-1{1'b0}}, 1'b1};

////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//

assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);

// Guard Bit ...
always @(posedge clk or posedge rst)
	if(rst)						gb <= 1'b0;
	else
	if(clr)						gb <= 1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <= 1'b1;
	else
	if(re)						gb <= 1'b0;

endmodule

module dpram_512_40bit #(
	parameter DWIDTH = 40,
	parameter AWIDTH = 9
  )
  (
	clk,
	address_a,
	address_b,
	wren_a,
	wren_b,
	data_a,
	data_b,
	out_a,
	out_b
);

parameter NUM_WORDS=1<<AWIDTH;

input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

	reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];

	always @ (posedge clk) begin
		if (wren_a) begin
			ram[address_a] <= data_a;
		end
		else begin
			out_a <= ram[address_a];
		end
	end
	  
	always @ (posedge clk) begin 
		if (wren_b) begin
			ram[address_b] <= data_b;
		end 
		else begin
			out_b <= ram[address_b];
		end
	end

`else
defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

	dual_port_ram u_dual_port_ram(
	.addr1(address_a),
	.we1(wren_a),
	.data1(data_a),
	.out1(out_a),
	.addr2(address_b),
	.we2(wren_b),
	.data2(data_b),
	.out2(out_b),
	.clk(clk)
	);

`endif

endmodule

module dsp_chain_3_int_sop_2 (clk,reset,ax1,ay1,bx1,by1,ax2,ay2,bx2,by2,ax3,ay3,bx3,by3,result);

input clk; 
input reset; 
input [17:0] ax1, bx1, ax2, bx2, ax3, bx3; 
input [18:0] ay1, by1, ay2, by2, ay3, by3; 
output reg [36:0] result; 

wire [36:0] chainout0, chainout1, chainout2; 
wire [36:0] chainin0, chainin1, chainin2; 
wire [36:0] resulta1, resulta2, resulta3;

assign chainin0 = 37'd0;

int_sop_2_dspchain inst1 (.clk(clk),.reset(reset),.ax(ax1),.bx(bx1),.ay(ay1),.by(by1),.mode_sigs(11'd0),.chainin(chainin0),.resulta(resulta1),.chainout(chainout0));
int_sop_2_dspchain inst2 (.clk(clk),.reset(reset),.ax(ax2),.bx(bx2),.ay(ay2),.by(by2),.mode_sigs(11'd0),.chainin(chainout0),.resulta(resulta2),.chainout(chainout1));
int_sop_2_dspchain inst3 (.clk(clk),.reset(reset),.ax(ax3),.bx(bx3),.ay(ay3),.by(by3),.mode_sigs(11'd0),.chainin(chainout1),.resulta(resulta3),.chainout(chainout2));

assign result = resulta3;


endmodule 
module dsp_chain_2_int_sop_2 (clk,reset,ax1,ay1,bx1,by1,ax2,ay2,bx2,by2,result);

input clk; 
input reset; 
input [17:0] ax1, bx1, ax2, bx2; 
input [18:0] ay1, by1, ay2, by2; 
output reg [36:0] result; 

wire [36:0] chainout0, chainout1; 
wire [36:0] chainin0, chainin1; 
wire [36:0] resulta1, resulta2;

assign chainin0 = 37'd0;

int_sop_2_dspchain inst1 (.clk(clk),.reset(reset),.ax(ax1),.bx(bx1),.ay(ay1),.by(by1),.mode_sigs(11'd0),.chainin(chainin0),.resulta(resulta1),.chainout(chainout0));
int_sop_2_dspchain inst2 (.clk(clk),.reset(reset),.ax(ax2),.bx(bx2),.ay(ay2),.by(by2),.mode_sigs(11'd0),.chainin(chainout0),.resulta(resulta2),.chainout(chainout1));

assign result = resulta2;


endmodule 
