
module top (input clk, input reset,input [729:0] top_inp, output [303:0] top_outp); 
 


 wire [207:0] inp_spram1;
wire [159:0] outp_spram1;

spram_2048_40bit_module_4 spram1 (.clk(clk),.reset(reset),.inp(inp_spram1),.outp(outp_spram1)); 


 wire [794:0] inp_dot1;
wire [815:0] outp_dot1;

tensor_block_bf16_module_3 dot1 (.clk(clk),.reset(reset),.inp(inp_dot1),.outp(outp_dot1)); 
wire [159:0] inp_interface_1; 
wire [794:0] outp_interface_1; 

interface_1 inst_interface_1(.clk(clk),.reset(reset),.inp(inp_interface_1),.outp(outp_interface_1)); 


 wire [417:0] inp_sys_array1;
wire [223:0] outp_sys_array1;

systolic_array_4_fp16bit_1 sys_array1 (.clk(clk),.reset(reset),.inp(inp_sys_array1),.outp(outp_sys_array1)); 
wire [351:0] inp_interface_2; 
wire [417:0] outp_interface_2; 

interface_2 inst_interface_2(.clk(clk),.reset(reset),.inp(inp_interface_2),.outp(outp_interface_2)); 


 wire [835:0] inp_sys_array2;
wire [447:0] outp_sys_array2;

systolic_array_4_fp16bit_2 sys_array2 (.clk(clk),.reset(reset),.inp(inp_sys_array2),.outp(outp_sys_array2)); 
wire [815:0] inp_interface_3; 
wire [835:0] outp_interface_3; 

interface_3 inst_interface_3(.clk(clk),.reset(reset),.inp(inp_interface_3),.outp(outp_interface_3)); 


 wire [835:0] inp_sys_array3;
wire [447:0] outp_sys_array3;

systolic_array_4_fp16bit_2 sys_array3 (.clk(clk),.reset(reset),.inp(inp_sys_array3),.outp(outp_sys_array3)); 
wire [815:0] inp_interface_4; 
wire [835:0] outp_interface_4; 

interface_4 inst_interface_4(.clk(clk),.reset(reset),.inp(inp_interface_4),.outp(outp_interface_4)); 


 wire [875:0] inp_spram2;
wire [719:0] outp_spram2;

spram_4096_60bit_module_12 spram2 (.clk(clk),.reset(reset),.inp(inp_spram2),.outp(outp_spram2)); 
wire [223:0] inp_interface_5; 
wire [875:0] outp_interface_5; 

interface_5 inst_interface_5(.clk(clk),.reset(reset),.inp(inp_interface_5),.outp(outp_interface_5)); 


 wire [1535:0] inp_adder_tree1;
wire [191:0] outp_adder_tree1;

adder_tree_4_8bit_12 adder_tree1 (.clk(clk),.reset(reset),.inp(inp_adder_tree1),.outp(outp_adder_tree1)); 
wire [4015:0] inp_interface_6; 
wire [1535:0] outp_interface_6; 

interface_6 inst_interface_6(.clk(clk),.reset(reset),.inp(inp_interface_6),.outp(outp_interface_6)); 


 wire [3179:0] inp_spram3;
wire [2399:0] outp_spram3;

spram_4096_40bit_module_60 spram3 (.clk(clk),.reset(reset),.inp(inp_spram3),.outp(outp_spram3)); 
wire [1663:0] inp_interface_7; 
wire [3179:0] outp_interface_7; 

interface_7 inst_interface_7(.clk(clk),.reset(reset),.inp(inp_interface_7),.outp(outp_interface_7)); 


 wire [529:0] inp_dot2;
wire [543:0] outp_dot2;

tensor_block_bf16_module_2 dot2 (.clk(clk),.reset(reset),.inp(inp_dot2),.outp(outp_dot2)); 
wire [191:0] inp_interface_8; 
wire [529:0] outp_interface_8; 

interface_8 inst_interface_8(.clk(clk),.reset(reset),.inp(inp_interface_8),.outp(outp_interface_8)); 


 wire [417:0] inp_sys_array4;
wire [223:0] outp_sys_array4;

systolic_array_4_fp16bit_1 sys_array4 (.clk(clk),.reset(reset),.inp(inp_sys_array4),.outp(outp_sys_array4)); 


 wire [1055:0] inp_adder_tree2;
wire [127:0] outp_adder_tree2;

adder_tree_3_fp16bit_8 adder_tree2 (.clk(clk),.reset(reset),.inp(inp_adder_tree2),.outp(outp_adder_tree2)); 
wire [2623:0] inp_interface_10; 
wire [1055:0] outp_interface_10; 

interface_10 inst_interface_10(.clk(clk),.reset(reset),.inp(inp_interface_10),.outp(outp_interface_10)); 


 wire [103:0] inp_spram4;
wire [79:0] outp_spram4;

spram_2048_40bit_module_2 spram4 (.clk(clk),.reset(reset),.inp(inp_spram4),.outp(outp_spram4)); 


 wire [511:0] inp_adder_tree3;
wire [127:0] outp_adder_tree3;

adder_tree_3_16bit_4 adder_tree3 (.clk(clk),.reset(reset),.inp(inp_adder_tree3),.outp(outp_adder_tree3)); 
wire [303:0] inp_interface_12; 
wire [511:0] outp_interface_12; 

interface_12 inst_interface_12(.clk(clk),.reset(reset),.inp(inp_interface_12),.outp(outp_interface_12)); 


 wire [1319:0] inp_adder_tree4;
wire [159:0] outp_adder_tree4;

adder_tree_3_fp16bit_10 adder_tree4 (.clk(clk),.reset(reset),.inp(inp_adder_tree4),.outp(outp_adder_tree4)); 
wire [4143:0] inp_interface_13; 
wire [1319:0] outp_interface_13; 

interface_13 inst_interface_13(.clk(clk),.reset(reset),.inp(inp_interface_13),.outp(outp_interface_13)); 


 wire [1055:0] inp_adder_tree5;
wire [127:0] outp_adder_tree5;

adder_tree_3_fp16bit_8 adder_tree5 (.clk(clk),.reset(reset),.inp(inp_adder_tree5),.outp(outp_adder_tree5)); 
wire [2687:0] inp_interface_14; 
wire [1055:0] outp_interface_14; 

interface_14 inst_interface_14(.clk(clk),.reset(reset),.inp(inp_interface_14),.outp(outp_interface_14)); 


 wire [1253:0] inp_sys_array5;
wire [671:0] outp_sys_array5;

systolic_array_4_fp16bit_3 sys_array5 (.clk(clk),.reset(reset),.inp(inp_sys_array5),.outp(outp_sys_array5)); 
wire [975:0] inp_interface_15; 
wire [1253:0] outp_interface_15; 

interface_15 inst_interface_15(.clk(clk),.reset(reset),.inp(inp_interface_15),.outp(outp_interface_15)); 


 wire [417:0] inp_sys_array6;
wire [223:0] outp_sys_array6;

systolic_array_4_fp16bit_1 sys_array6 (.clk(clk),.reset(reset),.inp(inp_sys_array6),.outp(outp_sys_array6)); 
wire [127:0] inp_interface_16; 
wire [417:0] outp_interface_16; 

interface_16 inst_interface_16(.clk(clk),.reset(reset),.inp(inp_interface_16),.outp(outp_interface_16)); 


 wire [1271:0] inp_spram5;
wire [959:0] outp_spram5;

spram_4096_40bit_module_24 spram5 (.clk(clk),.reset(reset),.inp(inp_spram5),.outp(outp_spram5)); 
wire [287:0] inp_interface_17; 
wire [1271:0] outp_interface_17; 

interface_17 inst_interface_17(.clk(clk),.reset(reset),.inp(inp_interface_17),.outp(outp_interface_17)); 


 wire [794:0] inp_dot3;
wire [815:0] outp_dot3;

tensor_block_bf16_module_3 dot3 (.clk(clk),.reset(reset),.inp(inp_dot3),.outp(outp_dot3)); 
wire [959:0] inp_interface_18; 
wire [794:0] outp_interface_18; 

interface_18 inst_interface_18(.clk(clk),.reset(reset),.inp(inp_interface_18),.outp(outp_interface_18)); 


 wire [103:0] inp_spram6;
wire [79:0] outp_spram6;

spram_2048_40bit_module_2 spram6 (.clk(clk),.reset(reset),.inp(inp_spram6),.outp(outp_spram6)); 
wire [815:0] inp_interface_19; 
wire [103:0] outp_interface_19; 

interface_19 inst_interface_19(.clk(clk),.reset(reset),.inp(inp_interface_19),.outp(outp_interface_19)); 

assign inp_spram1 = top_inp[207:0]; 

assign inp_dot1 = outp_interface_1; 
assign inp_interface_1 = {outp_spram1}; 
 

assign inp_sys_array1 = outp_interface_2; 
assign inp_interface_2 = {outp_spram1,outp_adder_tree1}; 
 

assign inp_sys_array2 = outp_interface_3; 
assign inp_interface_3 = {outp_dot1}; 
 

assign inp_sys_array3 = outp_interface_4; 
assign inp_interface_4 = {outp_dot1}; 
 

assign inp_spram2 = outp_interface_5; 
assign inp_interface_5 = {outp_sys_array1}; 
 

assign inp_adder_tree1 = outp_interface_6; 
assign inp_interface_6 = {outp_spram2,outp_sys_array2,outp_sys_array3,outp_spram3}; 
 

assign inp_spram3 = outp_interface_7; 
assign inp_interface_7 = {outp_dot2,outp_sys_array3,outp_sys_array5}; 
 

assign inp_dot2 = outp_interface_8; 
assign inp_interface_8 = {outp_adder_tree1}; 
 

assign inp_sys_array4 = top_inp[625:208]; 

assign inp_adder_tree2 = outp_interface_10; 
assign inp_interface_10 = {outp_spram3,outp_sys_array4}; 
 

assign inp_spram4 = top_inp[729:626]; 

assign inp_adder_tree3 = outp_interface_12; 
assign inp_interface_12 = {outp_spram4,outp_sys_array4}; 
 

assign inp_adder_tree4 = outp_interface_13; 
assign inp_interface_13 = {outp_spram3,outp_sys_array5,outp_adder_tree2,outp_adder_tree3,outp_dot3}; 
 

assign inp_adder_tree5 = outp_interface_14; 
assign inp_interface_14 = {outp_spram3,outp_adder_tree4,outp_adder_tree3}; 
 

assign inp_sys_array5 = outp_interface_15; 
assign inp_interface_15 = {outp_spram1,outp_dot1}; 
 

assign inp_sys_array6 = outp_interface_16; 
assign top_outp[223:0] = outp_sys_array6; 
assign inp_interface_16 = {outp_adder_tree5}; 
 

assign inp_spram5 = outp_interface_17; 
assign inp_interface_17 = {outp_adder_tree4,outp_adder_tree5}; 
 

assign inp_dot3 = outp_interface_18; 
assign inp_interface_18 = {outp_spram5}; 
 

assign inp_spram6 = outp_interface_19; 
assign top_outp[303:224] = outp_spram6; 
assign inp_interface_19 = {outp_dot3}; 
 

 endmodule 


module interface_1(input [159:0] inp, output reg [794:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[159:0] <= inp ; 
outp[319:160] <= inp ; 
outp[479:320] <= inp ; 
outp[639:480] <= inp ; 
outp[794:640] <= inp[154:0] ; 
end 
endmodule 

module interface_2(input [351:0] inp, output reg [417:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[351:0] <= inp ; 
outp[417:352] <= inp[65:0] ; 
end 
endmodule 

module interface_3(input [815:0] inp, output reg [835:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[815:0] <= inp ; 
outp[835:816] <= inp[19:0] ; 
end 
endmodule 

module interface_4(input [815:0] inp, output reg [835:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[815:0] <= inp ; 
outp[835:816] <= inp[19:0] ; 
end 
endmodule 

module interface_5(input [223:0] inp, output reg [875:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[223:0] <= inp ; 
outp[447:224] <= inp ; 
outp[671:448] <= inp ; 
outp[875:672] <= inp[203:0] ; 
end 
endmodule 

module interface_6(input [4015:0] inp, output reg [1535:0] outp, input clk, input reset);
reg [4015:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [2007:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4015]),.i2(intermediate_reg_0[4014]),.o(intermediate_reg_1[2007]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4013]),.i2(intermediate_reg_0[4012]),.o(intermediate_reg_1[2006]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4011]),.i2(intermediate_reg_0[4010]),.o(intermediate_reg_1[2005]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4009]),.i2(intermediate_reg_0[4008]),.o(intermediate_reg_1[2004]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4007]),.i2(intermediate_reg_0[4006]),.o(intermediate_reg_1[2003]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4005]),.i2(intermediate_reg_0[4004]),.o(intermediate_reg_1[2002])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4003]),.i2(intermediate_reg_0[4002]),.o(intermediate_reg_1[2001]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4001]),.i2(intermediate_reg_0[4000]),.o(intermediate_reg_1[2000])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3999]),.i2(intermediate_reg_0[3998]),.o(intermediate_reg_1[1999]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3997]),.i2(intermediate_reg_0[3996]),.o(intermediate_reg_1[1998]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3995]),.i2(intermediate_reg_0[3994]),.o(intermediate_reg_1[1997])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3993]),.i2(intermediate_reg_0[3992]),.o(intermediate_reg_1[1996]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3991]),.i2(intermediate_reg_0[3990]),.o(intermediate_reg_1[1995])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3989]),.i2(intermediate_reg_0[3988]),.o(intermediate_reg_1[1994])); 
mux_module mux_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3987]),.i2(intermediate_reg_0[3986]),.o(intermediate_reg_1[1993]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3985]),.i2(intermediate_reg_0[3984]),.o(intermediate_reg_1[1992]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3983]),.i2(intermediate_reg_0[3982]),.o(intermediate_reg_1[1991])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3981]),.i2(intermediate_reg_0[3980]),.o(intermediate_reg_1[1990]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3979]),.i2(intermediate_reg_0[3978]),.o(intermediate_reg_1[1989]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3977]),.i2(intermediate_reg_0[3976]),.o(intermediate_reg_1[1988])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3975]),.i2(intermediate_reg_0[3974]),.o(intermediate_reg_1[1987])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3973]),.i2(intermediate_reg_0[3972]),.o(intermediate_reg_1[1986])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3971]),.i2(intermediate_reg_0[3970]),.o(intermediate_reg_1[1985]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3969]),.i2(intermediate_reg_0[3968]),.o(intermediate_reg_1[1984])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3967]),.i2(intermediate_reg_0[3966]),.o(intermediate_reg_1[1983]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3965]),.i2(intermediate_reg_0[3964]),.o(intermediate_reg_1[1982]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3963]),.i2(intermediate_reg_0[3962]),.o(intermediate_reg_1[1981]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3961]),.i2(intermediate_reg_0[3960]),.o(intermediate_reg_1[1980]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3959]),.i2(intermediate_reg_0[3958]),.o(intermediate_reg_1[1979]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3957]),.i2(intermediate_reg_0[3956]),.o(intermediate_reg_1[1978])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3955]),.i2(intermediate_reg_0[3954]),.o(intermediate_reg_1[1977]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3953]),.i2(intermediate_reg_0[3952]),.o(intermediate_reg_1[1976]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3951]),.i2(intermediate_reg_0[3950]),.o(intermediate_reg_1[1975]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3949]),.i2(intermediate_reg_0[3948]),.o(intermediate_reg_1[1974])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3947]),.i2(intermediate_reg_0[3946]),.o(intermediate_reg_1[1973]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3945]),.i2(intermediate_reg_0[3944]),.o(intermediate_reg_1[1972]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3943]),.i2(intermediate_reg_0[3942]),.o(intermediate_reg_1[1971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3941]),.i2(intermediate_reg_0[3940]),.o(intermediate_reg_1[1970]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3939]),.i2(intermediate_reg_0[3938]),.o(intermediate_reg_1[1969])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3937]),.i2(intermediate_reg_0[3936]),.o(intermediate_reg_1[1968]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3935]),.i2(intermediate_reg_0[3934]),.o(intermediate_reg_1[1967])); 
mux_module mux_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3933]),.i2(intermediate_reg_0[3932]),.o(intermediate_reg_1[1966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3931]),.i2(intermediate_reg_0[3930]),.o(intermediate_reg_1[1965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3929]),.i2(intermediate_reg_0[3928]),.o(intermediate_reg_1[1964]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3927]),.i2(intermediate_reg_0[3926]),.o(intermediate_reg_1[1963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3925]),.i2(intermediate_reg_0[3924]),.o(intermediate_reg_1[1962]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3923]),.i2(intermediate_reg_0[3922]),.o(intermediate_reg_1[1961])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3921]),.i2(intermediate_reg_0[3920]),.o(intermediate_reg_1[1960])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3919]),.i2(intermediate_reg_0[3918]),.o(intermediate_reg_1[1959])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3917]),.i2(intermediate_reg_0[3916]),.o(intermediate_reg_1[1958]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3915]),.i2(intermediate_reg_0[3914]),.o(intermediate_reg_1[1957]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3913]),.i2(intermediate_reg_0[3912]),.o(intermediate_reg_1[1956]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3911]),.i2(intermediate_reg_0[3910]),.o(intermediate_reg_1[1955])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3909]),.i2(intermediate_reg_0[3908]),.o(intermediate_reg_1[1954]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3907]),.i2(intermediate_reg_0[3906]),.o(intermediate_reg_1[1953]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3905]),.i2(intermediate_reg_0[3904]),.o(intermediate_reg_1[1952])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3903]),.i2(intermediate_reg_0[3902]),.o(intermediate_reg_1[1951])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3901]),.i2(intermediate_reg_0[3900]),.o(intermediate_reg_1[1950]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3899]),.i2(intermediate_reg_0[3898]),.o(intermediate_reg_1[1949])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3897]),.i2(intermediate_reg_0[3896]),.o(intermediate_reg_1[1948]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3895]),.i2(intermediate_reg_0[3894]),.o(intermediate_reg_1[1947])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3893]),.i2(intermediate_reg_0[3892]),.o(intermediate_reg_1[1946])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3891]),.i2(intermediate_reg_0[3890]),.o(intermediate_reg_1[1945]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3889]),.i2(intermediate_reg_0[3888]),.o(intermediate_reg_1[1944]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3887]),.i2(intermediate_reg_0[3886]),.o(intermediate_reg_1[1943])); 
mux_module mux_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3885]),.i2(intermediate_reg_0[3884]),.o(intermediate_reg_1[1942]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3883]),.i2(intermediate_reg_0[3882]),.o(intermediate_reg_1[1941]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3881]),.i2(intermediate_reg_0[3880]),.o(intermediate_reg_1[1940]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3879]),.i2(intermediate_reg_0[3878]),.o(intermediate_reg_1[1939])); 
mux_module mux_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3877]),.i2(intermediate_reg_0[3876]),.o(intermediate_reg_1[1938]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3875]),.i2(intermediate_reg_0[3874]),.o(intermediate_reg_1[1937])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3873]),.i2(intermediate_reg_0[3872]),.o(intermediate_reg_1[1936]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3871]),.i2(intermediate_reg_0[3870]),.o(intermediate_reg_1[1935]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3869]),.i2(intermediate_reg_0[3868]),.o(intermediate_reg_1[1934]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3867]),.i2(intermediate_reg_0[3866]),.o(intermediate_reg_1[1933])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3865]),.i2(intermediate_reg_0[3864]),.o(intermediate_reg_1[1932]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3863]),.i2(intermediate_reg_0[3862]),.o(intermediate_reg_1[1931]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3861]),.i2(intermediate_reg_0[3860]),.o(intermediate_reg_1[1930]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3859]),.i2(intermediate_reg_0[3858]),.o(intermediate_reg_1[1929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3857]),.i2(intermediate_reg_0[3856]),.o(intermediate_reg_1[1928]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3855]),.i2(intermediate_reg_0[3854]),.o(intermediate_reg_1[1927])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3853]),.i2(intermediate_reg_0[3852]),.o(intermediate_reg_1[1926])); 
xor_module xor_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3851]),.i2(intermediate_reg_0[3850]),.o(intermediate_reg_1[1925])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3849]),.i2(intermediate_reg_0[3848]),.o(intermediate_reg_1[1924])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3847]),.i2(intermediate_reg_0[3846]),.o(intermediate_reg_1[1923])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3845]),.i2(intermediate_reg_0[3844]),.o(intermediate_reg_1[1922]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3843]),.i2(intermediate_reg_0[3842]),.o(intermediate_reg_1[1921])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3841]),.i2(intermediate_reg_0[3840]),.o(intermediate_reg_1[1920])); 
mux_module mux_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3839]),.i2(intermediate_reg_0[3838]),.o(intermediate_reg_1[1919]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3837]),.i2(intermediate_reg_0[3836]),.o(intermediate_reg_1[1918])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3835]),.i2(intermediate_reg_0[3834]),.o(intermediate_reg_1[1917])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3833]),.i2(intermediate_reg_0[3832]),.o(intermediate_reg_1[1916])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3831]),.i2(intermediate_reg_0[3830]),.o(intermediate_reg_1[1915])); 
mux_module mux_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3829]),.i2(intermediate_reg_0[3828]),.o(intermediate_reg_1[1914]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3827]),.i2(intermediate_reg_0[3826]),.o(intermediate_reg_1[1913]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3825]),.i2(intermediate_reg_0[3824]),.o(intermediate_reg_1[1912]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3823]),.i2(intermediate_reg_0[3822]),.o(intermediate_reg_1[1911]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3821]),.i2(intermediate_reg_0[3820]),.o(intermediate_reg_1[1910])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3819]),.i2(intermediate_reg_0[3818]),.o(intermediate_reg_1[1909])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3817]),.i2(intermediate_reg_0[3816]),.o(intermediate_reg_1[1908])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3815]),.i2(intermediate_reg_0[3814]),.o(intermediate_reg_1[1907])); 
mux_module mux_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3813]),.i2(intermediate_reg_0[3812]),.o(intermediate_reg_1[1906]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3811]),.i2(intermediate_reg_0[3810]),.o(intermediate_reg_1[1905])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3809]),.i2(intermediate_reg_0[3808]),.o(intermediate_reg_1[1904]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3807]),.i2(intermediate_reg_0[3806]),.o(intermediate_reg_1[1903]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3805]),.i2(intermediate_reg_0[3804]),.o(intermediate_reg_1[1902])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3803]),.i2(intermediate_reg_0[3802]),.o(intermediate_reg_1[1901])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3801]),.i2(intermediate_reg_0[3800]),.o(intermediate_reg_1[1900]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3799]),.i2(intermediate_reg_0[3798]),.o(intermediate_reg_1[1899])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3797]),.i2(intermediate_reg_0[3796]),.o(intermediate_reg_1[1898])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3795]),.i2(intermediate_reg_0[3794]),.o(intermediate_reg_1[1897])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3793]),.i2(intermediate_reg_0[3792]),.o(intermediate_reg_1[1896]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3791]),.i2(intermediate_reg_0[3790]),.o(intermediate_reg_1[1895]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3789]),.i2(intermediate_reg_0[3788]),.o(intermediate_reg_1[1894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3787]),.i2(intermediate_reg_0[3786]),.o(intermediate_reg_1[1893]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3785]),.i2(intermediate_reg_0[3784]),.o(intermediate_reg_1[1892])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3783]),.i2(intermediate_reg_0[3782]),.o(intermediate_reg_1[1891]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3781]),.i2(intermediate_reg_0[3780]),.o(intermediate_reg_1[1890])); 
mux_module mux_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3779]),.i2(intermediate_reg_0[3778]),.o(intermediate_reg_1[1889]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3777]),.i2(intermediate_reg_0[3776]),.o(intermediate_reg_1[1888]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3775]),.i2(intermediate_reg_0[3774]),.o(intermediate_reg_1[1887])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3773]),.i2(intermediate_reg_0[3772]),.o(intermediate_reg_1[1886]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3771]),.i2(intermediate_reg_0[3770]),.o(intermediate_reg_1[1885]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3769]),.i2(intermediate_reg_0[3768]),.o(intermediate_reg_1[1884]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3767]),.i2(intermediate_reg_0[3766]),.o(intermediate_reg_1[1883])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3765]),.i2(intermediate_reg_0[3764]),.o(intermediate_reg_1[1882])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3763]),.i2(intermediate_reg_0[3762]),.o(intermediate_reg_1[1881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3761]),.i2(intermediate_reg_0[3760]),.o(intermediate_reg_1[1880]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3759]),.i2(intermediate_reg_0[3758]),.o(intermediate_reg_1[1879]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3757]),.i2(intermediate_reg_0[3756]),.o(intermediate_reg_1[1878])); 
xor_module xor_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3755]),.i2(intermediate_reg_0[3754]),.o(intermediate_reg_1[1877])); 
mux_module mux_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3753]),.i2(intermediate_reg_0[3752]),.o(intermediate_reg_1[1876]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3751]),.i2(intermediate_reg_0[3750]),.o(intermediate_reg_1[1875])); 
mux_module mux_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3749]),.i2(intermediate_reg_0[3748]),.o(intermediate_reg_1[1874]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3747]),.i2(intermediate_reg_0[3746]),.o(intermediate_reg_1[1873]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3745]),.i2(intermediate_reg_0[3744]),.o(intermediate_reg_1[1872]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3743]),.i2(intermediate_reg_0[3742]),.o(intermediate_reg_1[1871])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3741]),.i2(intermediate_reg_0[3740]),.o(intermediate_reg_1[1870]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3739]),.i2(intermediate_reg_0[3738]),.o(intermediate_reg_1[1869])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3737]),.i2(intermediate_reg_0[3736]),.o(intermediate_reg_1[1868])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3735]),.i2(intermediate_reg_0[3734]),.o(intermediate_reg_1[1867])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3733]),.i2(intermediate_reg_0[3732]),.o(intermediate_reg_1[1866]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3731]),.i2(intermediate_reg_0[3730]),.o(intermediate_reg_1[1865])); 
mux_module mux_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3729]),.i2(intermediate_reg_0[3728]),.o(intermediate_reg_1[1864]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3727]),.i2(intermediate_reg_0[3726]),.o(intermediate_reg_1[1863])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3725]),.i2(intermediate_reg_0[3724]),.o(intermediate_reg_1[1862]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3723]),.i2(intermediate_reg_0[3722]),.o(intermediate_reg_1[1861])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3721]),.i2(intermediate_reg_0[3720]),.o(intermediate_reg_1[1860])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3719]),.i2(intermediate_reg_0[3718]),.o(intermediate_reg_1[1859]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3717]),.i2(intermediate_reg_0[3716]),.o(intermediate_reg_1[1858]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3715]),.i2(intermediate_reg_0[3714]),.o(intermediate_reg_1[1857])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3713]),.i2(intermediate_reg_0[3712]),.o(intermediate_reg_1[1856])); 
mux_module mux_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3711]),.i2(intermediate_reg_0[3710]),.o(intermediate_reg_1[1855]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3709]),.i2(intermediate_reg_0[3708]),.o(intermediate_reg_1[1854])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3707]),.i2(intermediate_reg_0[3706]),.o(intermediate_reg_1[1853])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3705]),.i2(intermediate_reg_0[3704]),.o(intermediate_reg_1[1852])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3703]),.i2(intermediate_reg_0[3702]),.o(intermediate_reg_1[1851])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3701]),.i2(intermediate_reg_0[3700]),.o(intermediate_reg_1[1850])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3699]),.i2(intermediate_reg_0[3698]),.o(intermediate_reg_1[1849])); 
mux_module mux_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3697]),.i2(intermediate_reg_0[3696]),.o(intermediate_reg_1[1848]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3695]),.i2(intermediate_reg_0[3694]),.o(intermediate_reg_1[1847]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3693]),.i2(intermediate_reg_0[3692]),.o(intermediate_reg_1[1846])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3691]),.i2(intermediate_reg_0[3690]),.o(intermediate_reg_1[1845]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3689]),.i2(intermediate_reg_0[3688]),.o(intermediate_reg_1[1844]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3687]),.i2(intermediate_reg_0[3686]),.o(intermediate_reg_1[1843])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3685]),.i2(intermediate_reg_0[3684]),.o(intermediate_reg_1[1842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3683]),.i2(intermediate_reg_0[3682]),.o(intermediate_reg_1[1841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3681]),.i2(intermediate_reg_0[3680]),.o(intermediate_reg_1[1840]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3679]),.i2(intermediate_reg_0[3678]),.o(intermediate_reg_1[1839]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3677]),.i2(intermediate_reg_0[3676]),.o(intermediate_reg_1[1838])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3675]),.i2(intermediate_reg_0[3674]),.o(intermediate_reg_1[1837])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3673]),.i2(intermediate_reg_0[3672]),.o(intermediate_reg_1[1836])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3671]),.i2(intermediate_reg_0[3670]),.o(intermediate_reg_1[1835]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3669]),.i2(intermediate_reg_0[3668]),.o(intermediate_reg_1[1834])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3667]),.i2(intermediate_reg_0[3666]),.o(intermediate_reg_1[1833])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3665]),.i2(intermediate_reg_0[3664]),.o(intermediate_reg_1[1832]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3663]),.i2(intermediate_reg_0[3662]),.o(intermediate_reg_1[1831])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3661]),.i2(intermediate_reg_0[3660]),.o(intermediate_reg_1[1830]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3659]),.i2(intermediate_reg_0[3658]),.o(intermediate_reg_1[1829])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3657]),.i2(intermediate_reg_0[3656]),.o(intermediate_reg_1[1828])); 
mux_module mux_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3655]),.i2(intermediate_reg_0[3654]),.o(intermediate_reg_1[1827]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3653]),.i2(intermediate_reg_0[3652]),.o(intermediate_reg_1[1826])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3651]),.i2(intermediate_reg_0[3650]),.o(intermediate_reg_1[1825])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3649]),.i2(intermediate_reg_0[3648]),.o(intermediate_reg_1[1824]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3647]),.i2(intermediate_reg_0[3646]),.o(intermediate_reg_1[1823])); 
xor_module xor_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3645]),.i2(intermediate_reg_0[3644]),.o(intermediate_reg_1[1822])); 
xor_module xor_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3643]),.i2(intermediate_reg_0[3642]),.o(intermediate_reg_1[1821])); 
xor_module xor_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3641]),.i2(intermediate_reg_0[3640]),.o(intermediate_reg_1[1820])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3639]),.i2(intermediate_reg_0[3638]),.o(intermediate_reg_1[1819])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3637]),.i2(intermediate_reg_0[3636]),.o(intermediate_reg_1[1818]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3635]),.i2(intermediate_reg_0[3634]),.o(intermediate_reg_1[1817]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3633]),.i2(intermediate_reg_0[3632]),.o(intermediate_reg_1[1816])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3631]),.i2(intermediate_reg_0[3630]),.o(intermediate_reg_1[1815]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3629]),.i2(intermediate_reg_0[3628]),.o(intermediate_reg_1[1814])); 
xor_module xor_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3627]),.i2(intermediate_reg_0[3626]),.o(intermediate_reg_1[1813])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3625]),.i2(intermediate_reg_0[3624]),.o(intermediate_reg_1[1812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3623]),.i2(intermediate_reg_0[3622]),.o(intermediate_reg_1[1811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3621]),.i2(intermediate_reg_0[3620]),.o(intermediate_reg_1[1810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3619]),.i2(intermediate_reg_0[3618]),.o(intermediate_reg_1[1809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3617]),.i2(intermediate_reg_0[3616]),.o(intermediate_reg_1[1808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3615]),.i2(intermediate_reg_0[3614]),.o(intermediate_reg_1[1807]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3613]),.i2(intermediate_reg_0[3612]),.o(intermediate_reg_1[1806]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3611]),.i2(intermediate_reg_0[3610]),.o(intermediate_reg_1[1805])); 
xor_module xor_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3609]),.i2(intermediate_reg_0[3608]),.o(intermediate_reg_1[1804])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3607]),.i2(intermediate_reg_0[3606]),.o(intermediate_reg_1[1803]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3605]),.i2(intermediate_reg_0[3604]),.o(intermediate_reg_1[1802])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3603]),.i2(intermediate_reg_0[3602]),.o(intermediate_reg_1[1801]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3601]),.i2(intermediate_reg_0[3600]),.o(intermediate_reg_1[1800])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3599]),.i2(intermediate_reg_0[3598]),.o(intermediate_reg_1[1799]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3597]),.i2(intermediate_reg_0[3596]),.o(intermediate_reg_1[1798])); 
xor_module xor_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3595]),.i2(intermediate_reg_0[3594]),.o(intermediate_reg_1[1797])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3593]),.i2(intermediate_reg_0[3592]),.o(intermediate_reg_1[1796])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3591]),.i2(intermediate_reg_0[3590]),.o(intermediate_reg_1[1795])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3589]),.i2(intermediate_reg_0[3588]),.o(intermediate_reg_1[1794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3587]),.i2(intermediate_reg_0[3586]),.o(intermediate_reg_1[1793]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3585]),.i2(intermediate_reg_0[3584]),.o(intermediate_reg_1[1792])); 
mux_module mux_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3583]),.i2(intermediate_reg_0[3582]),.o(intermediate_reg_1[1791]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3581]),.i2(intermediate_reg_0[3580]),.o(intermediate_reg_1[1790])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3579]),.i2(intermediate_reg_0[3578]),.o(intermediate_reg_1[1789]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3577]),.i2(intermediate_reg_0[3576]),.o(intermediate_reg_1[1788])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3575]),.i2(intermediate_reg_0[3574]),.o(intermediate_reg_1[1787])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3573]),.i2(intermediate_reg_0[3572]),.o(intermediate_reg_1[1786]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3571]),.i2(intermediate_reg_0[3570]),.o(intermediate_reg_1[1785])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3569]),.i2(intermediate_reg_0[3568]),.o(intermediate_reg_1[1784])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3567]),.i2(intermediate_reg_0[3566]),.o(intermediate_reg_1[1783])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3565]),.i2(intermediate_reg_0[3564]),.o(intermediate_reg_1[1782]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3563]),.i2(intermediate_reg_0[3562]),.o(intermediate_reg_1[1781])); 
mux_module mux_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3561]),.i2(intermediate_reg_0[3560]),.o(intermediate_reg_1[1780]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3559]),.i2(intermediate_reg_0[3558]),.o(intermediate_reg_1[1779])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3557]),.i2(intermediate_reg_0[3556]),.o(intermediate_reg_1[1778]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3555]),.i2(intermediate_reg_0[3554]),.o(intermediate_reg_1[1777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3553]),.i2(intermediate_reg_0[3552]),.o(intermediate_reg_1[1776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3551]),.i2(intermediate_reg_0[3550]),.o(intermediate_reg_1[1775]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3549]),.i2(intermediate_reg_0[3548]),.o(intermediate_reg_1[1774])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3547]),.i2(intermediate_reg_0[3546]),.o(intermediate_reg_1[1773])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3545]),.i2(intermediate_reg_0[3544]),.o(intermediate_reg_1[1772]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3543]),.i2(intermediate_reg_0[3542]),.o(intermediate_reg_1[1771])); 
mux_module mux_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3541]),.i2(intermediate_reg_0[3540]),.o(intermediate_reg_1[1770]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3539]),.i2(intermediate_reg_0[3538]),.o(intermediate_reg_1[1769])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3537]),.i2(intermediate_reg_0[3536]),.o(intermediate_reg_1[1768]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3535]),.i2(intermediate_reg_0[3534]),.o(intermediate_reg_1[1767]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3533]),.i2(intermediate_reg_0[3532]),.o(intermediate_reg_1[1766]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3531]),.i2(intermediate_reg_0[3530]),.o(intermediate_reg_1[1765])); 
mux_module mux_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3529]),.i2(intermediate_reg_0[3528]),.o(intermediate_reg_1[1764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3527]),.i2(intermediate_reg_0[3526]),.o(intermediate_reg_1[1763]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3525]),.i2(intermediate_reg_0[3524]),.o(intermediate_reg_1[1762])); 
xor_module xor_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3523]),.i2(intermediate_reg_0[3522]),.o(intermediate_reg_1[1761])); 
mux_module mux_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3521]),.i2(intermediate_reg_0[3520]),.o(intermediate_reg_1[1760]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3519]),.i2(intermediate_reg_0[3518]),.o(intermediate_reg_1[1759])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3517]),.i2(intermediate_reg_0[3516]),.o(intermediate_reg_1[1758]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3515]),.i2(intermediate_reg_0[3514]),.o(intermediate_reg_1[1757])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3513]),.i2(intermediate_reg_0[3512]),.o(intermediate_reg_1[1756])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3511]),.i2(intermediate_reg_0[3510]),.o(intermediate_reg_1[1755]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3509]),.i2(intermediate_reg_0[3508]),.o(intermediate_reg_1[1754]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3507]),.i2(intermediate_reg_0[3506]),.o(intermediate_reg_1[1753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3505]),.i2(intermediate_reg_0[3504]),.o(intermediate_reg_1[1752]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3503]),.i2(intermediate_reg_0[3502]),.o(intermediate_reg_1[1751])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3501]),.i2(intermediate_reg_0[3500]),.o(intermediate_reg_1[1750])); 
mux_module mux_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3499]),.i2(intermediate_reg_0[3498]),.o(intermediate_reg_1[1749]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3497]),.i2(intermediate_reg_0[3496]),.o(intermediate_reg_1[1748])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3495]),.i2(intermediate_reg_0[3494]),.o(intermediate_reg_1[1747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3493]),.i2(intermediate_reg_0[3492]),.o(intermediate_reg_1[1746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3491]),.i2(intermediate_reg_0[3490]),.o(intermediate_reg_1[1745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3489]),.i2(intermediate_reg_0[3488]),.o(intermediate_reg_1[1744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3487]),.i2(intermediate_reg_0[3486]),.o(intermediate_reg_1[1743]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3485]),.i2(intermediate_reg_0[3484]),.o(intermediate_reg_1[1742]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3483]),.i2(intermediate_reg_0[3482]),.o(intermediate_reg_1[1741])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3481]),.i2(intermediate_reg_0[3480]),.o(intermediate_reg_1[1740])); 
mux_module mux_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3479]),.i2(intermediate_reg_0[3478]),.o(intermediate_reg_1[1739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3477]),.i2(intermediate_reg_0[3476]),.o(intermediate_reg_1[1738]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3475]),.i2(intermediate_reg_0[3474]),.o(intermediate_reg_1[1737])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3473]),.i2(intermediate_reg_0[3472]),.o(intermediate_reg_1[1736])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3471]),.i2(intermediate_reg_0[3470]),.o(intermediate_reg_1[1735]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3469]),.i2(intermediate_reg_0[3468]),.o(intermediate_reg_1[1734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3467]),.i2(intermediate_reg_0[3466]),.o(intermediate_reg_1[1733]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3465]),.i2(intermediate_reg_0[3464]),.o(intermediate_reg_1[1732]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3463]),.i2(intermediate_reg_0[3462]),.o(intermediate_reg_1[1731])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3461]),.i2(intermediate_reg_0[3460]),.o(intermediate_reg_1[1730])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3459]),.i2(intermediate_reg_0[3458]),.o(intermediate_reg_1[1729]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3457]),.i2(intermediate_reg_0[3456]),.o(intermediate_reg_1[1728]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3455]),.i2(intermediate_reg_0[3454]),.o(intermediate_reg_1[1727]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3453]),.i2(intermediate_reg_0[3452]),.o(intermediate_reg_1[1726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3451]),.i2(intermediate_reg_0[3450]),.o(intermediate_reg_1[1725]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3449]),.i2(intermediate_reg_0[3448]),.o(intermediate_reg_1[1724])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3447]),.i2(intermediate_reg_0[3446]),.o(intermediate_reg_1[1723]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3445]),.i2(intermediate_reg_0[3444]),.o(intermediate_reg_1[1722])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3443]),.i2(intermediate_reg_0[3442]),.o(intermediate_reg_1[1721])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3441]),.i2(intermediate_reg_0[3440]),.o(intermediate_reg_1[1720]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3439]),.i2(intermediate_reg_0[3438]),.o(intermediate_reg_1[1719]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3437]),.i2(intermediate_reg_0[3436]),.o(intermediate_reg_1[1718])); 
mux_module mux_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3435]),.i2(intermediate_reg_0[3434]),.o(intermediate_reg_1[1717]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3433]),.i2(intermediate_reg_0[3432]),.o(intermediate_reg_1[1716])); 
xor_module xor_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3431]),.i2(intermediate_reg_0[3430]),.o(intermediate_reg_1[1715])); 
mux_module mux_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3429]),.i2(intermediate_reg_0[3428]),.o(intermediate_reg_1[1714]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3427]),.i2(intermediate_reg_0[3426]),.o(intermediate_reg_1[1713])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3425]),.i2(intermediate_reg_0[3424]),.o(intermediate_reg_1[1712])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3423]),.i2(intermediate_reg_0[3422]),.o(intermediate_reg_1[1711])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3421]),.i2(intermediate_reg_0[3420]),.o(intermediate_reg_1[1710])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3419]),.i2(intermediate_reg_0[3418]),.o(intermediate_reg_1[1709])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3417]),.i2(intermediate_reg_0[3416]),.o(intermediate_reg_1[1708])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3415]),.i2(intermediate_reg_0[3414]),.o(intermediate_reg_1[1707])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3413]),.i2(intermediate_reg_0[3412]),.o(intermediate_reg_1[1706]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3411]),.i2(intermediate_reg_0[3410]),.o(intermediate_reg_1[1705])); 
xor_module xor_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3409]),.i2(intermediate_reg_0[3408]),.o(intermediate_reg_1[1704])); 
mux_module mux_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3407]),.i2(intermediate_reg_0[3406]),.o(intermediate_reg_1[1703]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3405]),.i2(intermediate_reg_0[3404]),.o(intermediate_reg_1[1702])); 
mux_module mux_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3403]),.i2(intermediate_reg_0[3402]),.o(intermediate_reg_1[1701]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3401]),.i2(intermediate_reg_0[3400]),.o(intermediate_reg_1[1700])); 
mux_module mux_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3399]),.i2(intermediate_reg_0[3398]),.o(intermediate_reg_1[1699]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3397]),.i2(intermediate_reg_0[3396]),.o(intermediate_reg_1[1698])); 
mux_module mux_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3395]),.i2(intermediate_reg_0[3394]),.o(intermediate_reg_1[1697]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3393]),.i2(intermediate_reg_0[3392]),.o(intermediate_reg_1[1696])); 
mux_module mux_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3391]),.i2(intermediate_reg_0[3390]),.o(intermediate_reg_1[1695]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3389]),.i2(intermediate_reg_0[3388]),.o(intermediate_reg_1[1694])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3387]),.i2(intermediate_reg_0[3386]),.o(intermediate_reg_1[1693]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3385]),.i2(intermediate_reg_0[3384]),.o(intermediate_reg_1[1692])); 
mux_module mux_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3383]),.i2(intermediate_reg_0[3382]),.o(intermediate_reg_1[1691]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3381]),.i2(intermediate_reg_0[3380]),.o(intermediate_reg_1[1690])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3379]),.i2(intermediate_reg_0[3378]),.o(intermediate_reg_1[1689])); 
mux_module mux_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3377]),.i2(intermediate_reg_0[3376]),.o(intermediate_reg_1[1688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3375]),.i2(intermediate_reg_0[3374]),.o(intermediate_reg_1[1687]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3373]),.i2(intermediate_reg_0[3372]),.o(intermediate_reg_1[1686])); 
mux_module mux_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3371]),.i2(intermediate_reg_0[3370]),.o(intermediate_reg_1[1685]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3369]),.i2(intermediate_reg_0[3368]),.o(intermediate_reg_1[1684])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3367]),.i2(intermediate_reg_0[3366]),.o(intermediate_reg_1[1683])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3365]),.i2(intermediate_reg_0[3364]),.o(intermediate_reg_1[1682])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3363]),.i2(intermediate_reg_0[3362]),.o(intermediate_reg_1[1681]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3361]),.i2(intermediate_reg_0[3360]),.o(intermediate_reg_1[1680])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3359]),.i2(intermediate_reg_0[3358]),.o(intermediate_reg_1[1679])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3357]),.i2(intermediate_reg_0[3356]),.o(intermediate_reg_1[1678])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3355]),.i2(intermediate_reg_0[3354]),.o(intermediate_reg_1[1677]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3353]),.i2(intermediate_reg_0[3352]),.o(intermediate_reg_1[1676])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3351]),.i2(intermediate_reg_0[3350]),.o(intermediate_reg_1[1675])); 
xor_module xor_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3349]),.i2(intermediate_reg_0[3348]),.o(intermediate_reg_1[1674])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3347]),.i2(intermediate_reg_0[3346]),.o(intermediate_reg_1[1673])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3345]),.i2(intermediate_reg_0[3344]),.o(intermediate_reg_1[1672]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3343]),.i2(intermediate_reg_0[3342]),.o(intermediate_reg_1[1671])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3341]),.i2(intermediate_reg_0[3340]),.o(intermediate_reg_1[1670])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3339]),.i2(intermediate_reg_0[3338]),.o(intermediate_reg_1[1669])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3337]),.i2(intermediate_reg_0[3336]),.o(intermediate_reg_1[1668])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3335]),.i2(intermediate_reg_0[3334]),.o(intermediate_reg_1[1667]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3333]),.i2(intermediate_reg_0[3332]),.o(intermediate_reg_1[1666])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3331]),.i2(intermediate_reg_0[3330]),.o(intermediate_reg_1[1665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3329]),.i2(intermediate_reg_0[3328]),.o(intermediate_reg_1[1664]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3327]),.i2(intermediate_reg_0[3326]),.o(intermediate_reg_1[1663])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3325]),.i2(intermediate_reg_0[3324]),.o(intermediate_reg_1[1662])); 
mux_module mux_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3323]),.i2(intermediate_reg_0[3322]),.o(intermediate_reg_1[1661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3321]),.i2(intermediate_reg_0[3320]),.o(intermediate_reg_1[1660]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3319]),.i2(intermediate_reg_0[3318]),.o(intermediate_reg_1[1659]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3317]),.i2(intermediate_reg_0[3316]),.o(intermediate_reg_1[1658])); 
mux_module mux_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3315]),.i2(intermediate_reg_0[3314]),.o(intermediate_reg_1[1657]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3313]),.i2(intermediate_reg_0[3312]),.o(intermediate_reg_1[1656])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3311]),.i2(intermediate_reg_0[3310]),.o(intermediate_reg_1[1655]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3309]),.i2(intermediate_reg_0[3308]),.o(intermediate_reg_1[1654]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3307]),.i2(intermediate_reg_0[3306]),.o(intermediate_reg_1[1653])); 
xor_module xor_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3305]),.i2(intermediate_reg_0[3304]),.o(intermediate_reg_1[1652])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3303]),.i2(intermediate_reg_0[3302]),.o(intermediate_reg_1[1651])); 
xor_module xor_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3301]),.i2(intermediate_reg_0[3300]),.o(intermediate_reg_1[1650])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3299]),.i2(intermediate_reg_0[3298]),.o(intermediate_reg_1[1649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3297]),.i2(intermediate_reg_0[3296]),.o(intermediate_reg_1[1648]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3295]),.i2(intermediate_reg_0[3294]),.o(intermediate_reg_1[1647])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3293]),.i2(intermediate_reg_0[3292]),.o(intermediate_reg_1[1646])); 
mux_module mux_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3291]),.i2(intermediate_reg_0[3290]),.o(intermediate_reg_1[1645]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3289]),.i2(intermediate_reg_0[3288]),.o(intermediate_reg_1[1644])); 
mux_module mux_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3287]),.i2(intermediate_reg_0[3286]),.o(intermediate_reg_1[1643]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3285]),.i2(intermediate_reg_0[3284]),.o(intermediate_reg_1[1642])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3283]),.i2(intermediate_reg_0[3282]),.o(intermediate_reg_1[1641])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3281]),.i2(intermediate_reg_0[3280]),.o(intermediate_reg_1[1640])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3279]),.i2(intermediate_reg_0[3278]),.o(intermediate_reg_1[1639]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3277]),.i2(intermediate_reg_0[3276]),.o(intermediate_reg_1[1638])); 
mux_module mux_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3275]),.i2(intermediate_reg_0[3274]),.o(intermediate_reg_1[1637]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3273]),.i2(intermediate_reg_0[3272]),.o(intermediate_reg_1[1636]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3271]),.i2(intermediate_reg_0[3270]),.o(intermediate_reg_1[1635])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3269]),.i2(intermediate_reg_0[3268]),.o(intermediate_reg_1[1634]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3267]),.i2(intermediate_reg_0[3266]),.o(intermediate_reg_1[1633])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3265]),.i2(intermediate_reg_0[3264]),.o(intermediate_reg_1[1632])); 
mux_module mux_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3263]),.i2(intermediate_reg_0[3262]),.o(intermediate_reg_1[1631]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3261]),.i2(intermediate_reg_0[3260]),.o(intermediate_reg_1[1630]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3259]),.i2(intermediate_reg_0[3258]),.o(intermediate_reg_1[1629])); 
mux_module mux_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3257]),.i2(intermediate_reg_0[3256]),.o(intermediate_reg_1[1628]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3255]),.i2(intermediate_reg_0[3254]),.o(intermediate_reg_1[1627])); 
xor_module xor_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3253]),.i2(intermediate_reg_0[3252]),.o(intermediate_reg_1[1626])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3251]),.i2(intermediate_reg_0[3250]),.o(intermediate_reg_1[1625])); 
xor_module xor_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3249]),.i2(intermediate_reg_0[3248]),.o(intermediate_reg_1[1624])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3247]),.i2(intermediate_reg_0[3246]),.o(intermediate_reg_1[1623])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3245]),.i2(intermediate_reg_0[3244]),.o(intermediate_reg_1[1622]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3243]),.i2(intermediate_reg_0[3242]),.o(intermediate_reg_1[1621])); 
xor_module xor_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3241]),.i2(intermediate_reg_0[3240]),.o(intermediate_reg_1[1620])); 
mux_module mux_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3239]),.i2(intermediate_reg_0[3238]),.o(intermediate_reg_1[1619]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3237]),.i2(intermediate_reg_0[3236]),.o(intermediate_reg_1[1618])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3235]),.i2(intermediate_reg_0[3234]),.o(intermediate_reg_1[1617])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3233]),.i2(intermediate_reg_0[3232]),.o(intermediate_reg_1[1616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3231]),.i2(intermediate_reg_0[3230]),.o(intermediate_reg_1[1615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3229]),.i2(intermediate_reg_0[3228]),.o(intermediate_reg_1[1614]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3227]),.i2(intermediate_reg_0[3226]),.o(intermediate_reg_1[1613])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3225]),.i2(intermediate_reg_0[3224]),.o(intermediate_reg_1[1612]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3223]),.i2(intermediate_reg_0[3222]),.o(intermediate_reg_1[1611]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3221]),.i2(intermediate_reg_0[3220]),.o(intermediate_reg_1[1610])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3219]),.i2(intermediate_reg_0[3218]),.o(intermediate_reg_1[1609])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3217]),.i2(intermediate_reg_0[3216]),.o(intermediate_reg_1[1608])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3215]),.i2(intermediate_reg_0[3214]),.o(intermediate_reg_1[1607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3213]),.i2(intermediate_reg_0[3212]),.o(intermediate_reg_1[1606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3211]),.i2(intermediate_reg_0[3210]),.o(intermediate_reg_1[1605]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3209]),.i2(intermediate_reg_0[3208]),.o(intermediate_reg_1[1604])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3207]),.i2(intermediate_reg_0[3206]),.o(intermediate_reg_1[1603])); 
xor_module xor_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3205]),.i2(intermediate_reg_0[3204]),.o(intermediate_reg_1[1602])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3203]),.i2(intermediate_reg_0[3202]),.o(intermediate_reg_1[1601])); 
xor_module xor_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3201]),.i2(intermediate_reg_0[3200]),.o(intermediate_reg_1[1600])); 
mux_module mux_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3199]),.i2(intermediate_reg_0[3198]),.o(intermediate_reg_1[1599]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3197]),.i2(intermediate_reg_0[3196]),.o(intermediate_reg_1[1598]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3195]),.i2(intermediate_reg_0[3194]),.o(intermediate_reg_1[1597])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3193]),.i2(intermediate_reg_0[3192]),.o(intermediate_reg_1[1596])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3191]),.i2(intermediate_reg_0[3190]),.o(intermediate_reg_1[1595])); 
mux_module mux_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3189]),.i2(intermediate_reg_0[3188]),.o(intermediate_reg_1[1594]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3187]),.i2(intermediate_reg_0[3186]),.o(intermediate_reg_1[1593])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3185]),.i2(intermediate_reg_0[3184]),.o(intermediate_reg_1[1592])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3183]),.i2(intermediate_reg_0[3182]),.o(intermediate_reg_1[1591])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3181]),.i2(intermediate_reg_0[3180]),.o(intermediate_reg_1[1590]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3179]),.i2(intermediate_reg_0[3178]),.o(intermediate_reg_1[1589])); 
xor_module xor_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3177]),.i2(intermediate_reg_0[3176]),.o(intermediate_reg_1[1588])); 
mux_module mux_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3175]),.i2(intermediate_reg_0[3174]),.o(intermediate_reg_1[1587]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3173]),.i2(intermediate_reg_0[3172]),.o(intermediate_reg_1[1586])); 
xor_module xor_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3171]),.i2(intermediate_reg_0[3170]),.o(intermediate_reg_1[1585])); 
xor_module xor_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3169]),.i2(intermediate_reg_0[3168]),.o(intermediate_reg_1[1584])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3167]),.i2(intermediate_reg_0[3166]),.o(intermediate_reg_1[1583])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3165]),.i2(intermediate_reg_0[3164]),.o(intermediate_reg_1[1582])); 
mux_module mux_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3163]),.i2(intermediate_reg_0[3162]),.o(intermediate_reg_1[1581]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3161]),.i2(intermediate_reg_0[3160]),.o(intermediate_reg_1[1580])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3159]),.i2(intermediate_reg_0[3158]),.o(intermediate_reg_1[1579])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3157]),.i2(intermediate_reg_0[3156]),.o(intermediate_reg_1[1578]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3155]),.i2(intermediate_reg_0[3154]),.o(intermediate_reg_1[1577])); 
xor_module xor_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3153]),.i2(intermediate_reg_0[3152]),.o(intermediate_reg_1[1576])); 
xor_module xor_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3151]),.i2(intermediate_reg_0[3150]),.o(intermediate_reg_1[1575])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3149]),.i2(intermediate_reg_0[3148]),.o(intermediate_reg_1[1574]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3147]),.i2(intermediate_reg_0[3146]),.o(intermediate_reg_1[1573])); 
mux_module mux_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3145]),.i2(intermediate_reg_0[3144]),.o(intermediate_reg_1[1572]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3143]),.i2(intermediate_reg_0[3142]),.o(intermediate_reg_1[1571]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3141]),.i2(intermediate_reg_0[3140]),.o(intermediate_reg_1[1570]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3139]),.i2(intermediate_reg_0[3138]),.o(intermediate_reg_1[1569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3137]),.i2(intermediate_reg_0[3136]),.o(intermediate_reg_1[1568]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3135]),.i2(intermediate_reg_0[3134]),.o(intermediate_reg_1[1567])); 
mux_module mux_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3133]),.i2(intermediate_reg_0[3132]),.o(intermediate_reg_1[1566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3131]),.i2(intermediate_reg_0[3130]),.o(intermediate_reg_1[1565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3129]),.i2(intermediate_reg_0[3128]),.o(intermediate_reg_1[1564]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3127]),.i2(intermediate_reg_0[3126]),.o(intermediate_reg_1[1563])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3125]),.i2(intermediate_reg_0[3124]),.o(intermediate_reg_1[1562])); 
mux_module mux_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3123]),.i2(intermediate_reg_0[3122]),.o(intermediate_reg_1[1561]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3121]),.i2(intermediate_reg_0[3120]),.o(intermediate_reg_1[1560]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3119]),.i2(intermediate_reg_0[3118]),.o(intermediate_reg_1[1559])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3117]),.i2(intermediate_reg_0[3116]),.o(intermediate_reg_1[1558]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3115]),.i2(intermediate_reg_0[3114]),.o(intermediate_reg_1[1557]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3113]),.i2(intermediate_reg_0[3112]),.o(intermediate_reg_1[1556]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3111]),.i2(intermediate_reg_0[3110]),.o(intermediate_reg_1[1555])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3109]),.i2(intermediate_reg_0[3108]),.o(intermediate_reg_1[1554])); 
mux_module mux_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3107]),.i2(intermediate_reg_0[3106]),.o(intermediate_reg_1[1553]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3105]),.i2(intermediate_reg_0[3104]),.o(intermediate_reg_1[1552])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3103]),.i2(intermediate_reg_0[3102]),.o(intermediate_reg_1[1551])); 
mux_module mux_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3101]),.i2(intermediate_reg_0[3100]),.o(intermediate_reg_1[1550]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3099]),.i2(intermediate_reg_0[3098]),.o(intermediate_reg_1[1549])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3097]),.i2(intermediate_reg_0[3096]),.o(intermediate_reg_1[1548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3095]),.i2(intermediate_reg_0[3094]),.o(intermediate_reg_1[1547]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3093]),.i2(intermediate_reg_0[3092]),.o(intermediate_reg_1[1546])); 
mux_module mux_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3091]),.i2(intermediate_reg_0[3090]),.o(intermediate_reg_1[1545]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3089]),.i2(intermediate_reg_0[3088]),.o(intermediate_reg_1[1544])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3087]),.i2(intermediate_reg_0[3086]),.o(intermediate_reg_1[1543])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3085]),.i2(intermediate_reg_0[3084]),.o(intermediate_reg_1[1542])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3083]),.i2(intermediate_reg_0[3082]),.o(intermediate_reg_1[1541]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3081]),.i2(intermediate_reg_0[3080]),.o(intermediate_reg_1[1540])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3079]),.i2(intermediate_reg_0[3078]),.o(intermediate_reg_1[1539])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3077]),.i2(intermediate_reg_0[3076]),.o(intermediate_reg_1[1538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3075]),.i2(intermediate_reg_0[3074]),.o(intermediate_reg_1[1537]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3073]),.i2(intermediate_reg_0[3072]),.o(intermediate_reg_1[1536])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3071]),.i2(intermediate_reg_0[3070]),.o(intermediate_reg_1[1535])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3069]),.i2(intermediate_reg_0[3068]),.o(intermediate_reg_1[1534]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3067]),.i2(intermediate_reg_0[3066]),.o(intermediate_reg_1[1533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3065]),.i2(intermediate_reg_0[3064]),.o(intermediate_reg_1[1532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3063]),.i2(intermediate_reg_0[3062]),.o(intermediate_reg_1[1531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3061]),.i2(intermediate_reg_0[3060]),.o(intermediate_reg_1[1530]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3059]),.i2(intermediate_reg_0[3058]),.o(intermediate_reg_1[1529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3057]),.i2(intermediate_reg_0[3056]),.o(intermediate_reg_1[1528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3055]),.i2(intermediate_reg_0[3054]),.o(intermediate_reg_1[1527]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3053]),.i2(intermediate_reg_0[3052]),.o(intermediate_reg_1[1526])); 
xor_module xor_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3051]),.i2(intermediate_reg_0[3050]),.o(intermediate_reg_1[1525])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3049]),.i2(intermediate_reg_0[3048]),.o(intermediate_reg_1[1524])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3047]),.i2(intermediate_reg_0[3046]),.o(intermediate_reg_1[1523])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3045]),.i2(intermediate_reg_0[3044]),.o(intermediate_reg_1[1522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3043]),.i2(intermediate_reg_0[3042]),.o(intermediate_reg_1[1521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3041]),.i2(intermediate_reg_0[3040]),.o(intermediate_reg_1[1520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3039]),.i2(intermediate_reg_0[3038]),.o(intermediate_reg_1[1519]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3037]),.i2(intermediate_reg_0[3036]),.o(intermediate_reg_1[1518])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3035]),.i2(intermediate_reg_0[3034]),.o(intermediate_reg_1[1517]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3033]),.i2(intermediate_reg_0[3032]),.o(intermediate_reg_1[1516])); 
xor_module xor_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3031]),.i2(intermediate_reg_0[3030]),.o(intermediate_reg_1[1515])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3029]),.i2(intermediate_reg_0[3028]),.o(intermediate_reg_1[1514]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3027]),.i2(intermediate_reg_0[3026]),.o(intermediate_reg_1[1513])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3025]),.i2(intermediate_reg_0[3024]),.o(intermediate_reg_1[1512])); 
mux_module mux_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3023]),.i2(intermediate_reg_0[3022]),.o(intermediate_reg_1[1511]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3021]),.i2(intermediate_reg_0[3020]),.o(intermediate_reg_1[1510])); 
mux_module mux_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3019]),.i2(intermediate_reg_0[3018]),.o(intermediate_reg_1[1509]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3017]),.i2(intermediate_reg_0[3016]),.o(intermediate_reg_1[1508])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3015]),.i2(intermediate_reg_0[3014]),.o(intermediate_reg_1[1507])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3013]),.i2(intermediate_reg_0[3012]),.o(intermediate_reg_1[1506])); 
mux_module mux_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3011]),.i2(intermediate_reg_0[3010]),.o(intermediate_reg_1[1505]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3009]),.i2(intermediate_reg_0[3008]),.o(intermediate_reg_1[1504])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3007]),.i2(intermediate_reg_0[3006]),.o(intermediate_reg_1[1503])); 
mux_module mux_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3005]),.i2(intermediate_reg_0[3004]),.o(intermediate_reg_1[1502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3003]),.i2(intermediate_reg_0[3002]),.o(intermediate_reg_1[1501]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3001]),.i2(intermediate_reg_0[3000]),.o(intermediate_reg_1[1500])); 
mux_module mux_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2999]),.i2(intermediate_reg_0[2998]),.o(intermediate_reg_1[1499]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2997]),.i2(intermediate_reg_0[2996]),.o(intermediate_reg_1[1498])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2995]),.i2(intermediate_reg_0[2994]),.o(intermediate_reg_1[1497]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2993]),.i2(intermediate_reg_0[2992]),.o(intermediate_reg_1[1496]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2991]),.i2(intermediate_reg_0[2990]),.o(intermediate_reg_1[1495])); 
mux_module mux_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2989]),.i2(intermediate_reg_0[2988]),.o(intermediate_reg_1[1494]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2987]),.i2(intermediate_reg_0[2986]),.o(intermediate_reg_1[1493]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2985]),.i2(intermediate_reg_0[2984]),.o(intermediate_reg_1[1492])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2983]),.i2(intermediate_reg_0[2982]),.o(intermediate_reg_1[1491])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2981]),.i2(intermediate_reg_0[2980]),.o(intermediate_reg_1[1490])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2979]),.i2(intermediate_reg_0[2978]),.o(intermediate_reg_1[1489]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2977]),.i2(intermediate_reg_0[2976]),.o(intermediate_reg_1[1488]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2975]),.i2(intermediate_reg_0[2974]),.o(intermediate_reg_1[1487])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2973]),.i2(intermediate_reg_0[2972]),.o(intermediate_reg_1[1486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2971]),.i2(intermediate_reg_0[2970]),.o(intermediate_reg_1[1485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2969]),.i2(intermediate_reg_0[2968]),.o(intermediate_reg_1[1484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2967]),.i2(intermediate_reg_0[2966]),.o(intermediate_reg_1[1483]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2965]),.i2(intermediate_reg_0[2964]),.o(intermediate_reg_1[1482])); 
mux_module mux_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2963]),.i2(intermediate_reg_0[2962]),.o(intermediate_reg_1[1481]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2961]),.i2(intermediate_reg_0[2960]),.o(intermediate_reg_1[1480])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2959]),.i2(intermediate_reg_0[2958]),.o(intermediate_reg_1[1479]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2957]),.i2(intermediate_reg_0[2956]),.o(intermediate_reg_1[1478]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2955]),.i2(intermediate_reg_0[2954]),.o(intermediate_reg_1[1477])); 
mux_module mux_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2953]),.i2(intermediate_reg_0[2952]),.o(intermediate_reg_1[1476]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2951]),.i2(intermediate_reg_0[2950]),.o(intermediate_reg_1[1475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2949]),.i2(intermediate_reg_0[2948]),.o(intermediate_reg_1[1474]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2947]),.i2(intermediate_reg_0[2946]),.o(intermediate_reg_1[1473])); 
mux_module mux_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2945]),.i2(intermediate_reg_0[2944]),.o(intermediate_reg_1[1472]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2943]),.i2(intermediate_reg_0[2942]),.o(intermediate_reg_1[1471])); 
xor_module xor_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2941]),.i2(intermediate_reg_0[2940]),.o(intermediate_reg_1[1470])); 
xor_module xor_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2939]),.i2(intermediate_reg_0[2938]),.o(intermediate_reg_1[1469])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2937]),.i2(intermediate_reg_0[2936]),.o(intermediate_reg_1[1468]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2935]),.i2(intermediate_reg_0[2934]),.o(intermediate_reg_1[1467])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2933]),.i2(intermediate_reg_0[2932]),.o(intermediate_reg_1[1466])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2931]),.i2(intermediate_reg_0[2930]),.o(intermediate_reg_1[1465])); 
mux_module mux_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2929]),.i2(intermediate_reg_0[2928]),.o(intermediate_reg_1[1464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2927]),.i2(intermediate_reg_0[2926]),.o(intermediate_reg_1[1463]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2925]),.i2(intermediate_reg_0[2924]),.o(intermediate_reg_1[1462])); 
mux_module mux_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2923]),.i2(intermediate_reg_0[2922]),.o(intermediate_reg_1[1461]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2921]),.i2(intermediate_reg_0[2920]),.o(intermediate_reg_1[1460])); 
mux_module mux_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2919]),.i2(intermediate_reg_0[2918]),.o(intermediate_reg_1[1459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2917]),.i2(intermediate_reg_0[2916]),.o(intermediate_reg_1[1458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2915]),.i2(intermediate_reg_0[2914]),.o(intermediate_reg_1[1457])); 
xor_module xor_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2913]),.i2(intermediate_reg_0[2912]),.o(intermediate_reg_1[1456])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2911]),.i2(intermediate_reg_0[2910]),.o(intermediate_reg_1[1455])); 
mux_module mux_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2909]),.i2(intermediate_reg_0[2908]),.o(intermediate_reg_1[1454]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2907]),.i2(intermediate_reg_0[2906]),.o(intermediate_reg_1[1453])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2905]),.i2(intermediate_reg_0[2904]),.o(intermediate_reg_1[1452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2903]),.i2(intermediate_reg_0[2902]),.o(intermediate_reg_1[1451]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2901]),.i2(intermediate_reg_0[2900]),.o(intermediate_reg_1[1450]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2899]),.i2(intermediate_reg_0[2898]),.o(intermediate_reg_1[1449])); 
mux_module mux_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2897]),.i2(intermediate_reg_0[2896]),.o(intermediate_reg_1[1448]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2895]),.i2(intermediate_reg_0[2894]),.o(intermediate_reg_1[1447]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2893]),.i2(intermediate_reg_0[2892]),.o(intermediate_reg_1[1446])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2891]),.i2(intermediate_reg_0[2890]),.o(intermediate_reg_1[1445]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2889]),.i2(intermediate_reg_0[2888]),.o(intermediate_reg_1[1444])); 
xor_module xor_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2887]),.i2(intermediate_reg_0[2886]),.o(intermediate_reg_1[1443])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2885]),.i2(intermediate_reg_0[2884]),.o(intermediate_reg_1[1442])); 
xor_module xor_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2883]),.i2(intermediate_reg_0[2882]),.o(intermediate_reg_1[1441])); 
mux_module mux_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2881]),.i2(intermediate_reg_0[2880]),.o(intermediate_reg_1[1440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2879]),.i2(intermediate_reg_0[2878]),.o(intermediate_reg_1[1439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2877]),.i2(intermediate_reg_0[2876]),.o(intermediate_reg_1[1438]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2875]),.i2(intermediate_reg_0[2874]),.o(intermediate_reg_1[1437]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2873]),.i2(intermediate_reg_0[2872]),.o(intermediate_reg_1[1436]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2871]),.i2(intermediate_reg_0[2870]),.o(intermediate_reg_1[1435])); 
xor_module xor_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2869]),.i2(intermediate_reg_0[2868]),.o(intermediate_reg_1[1434])); 
mux_module mux_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2867]),.i2(intermediate_reg_0[2866]),.o(intermediate_reg_1[1433]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2865]),.i2(intermediate_reg_0[2864]),.o(intermediate_reg_1[1432])); 
mux_module mux_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2863]),.i2(intermediate_reg_0[2862]),.o(intermediate_reg_1[1431]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2861]),.i2(intermediate_reg_0[2860]),.o(intermediate_reg_1[1430])); 
mux_module mux_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2859]),.i2(intermediate_reg_0[2858]),.o(intermediate_reg_1[1429]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2857]),.i2(intermediate_reg_0[2856]),.o(intermediate_reg_1[1428])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2855]),.i2(intermediate_reg_0[2854]),.o(intermediate_reg_1[1427])); 
mux_module mux_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2853]),.i2(intermediate_reg_0[2852]),.o(intermediate_reg_1[1426]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2851]),.i2(intermediate_reg_0[2850]),.o(intermediate_reg_1[1425]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2849]),.i2(intermediate_reg_0[2848]),.o(intermediate_reg_1[1424])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2847]),.i2(intermediate_reg_0[2846]),.o(intermediate_reg_1[1423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2845]),.i2(intermediate_reg_0[2844]),.o(intermediate_reg_1[1422]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2843]),.i2(intermediate_reg_0[2842]),.o(intermediate_reg_1[1421]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2841]),.i2(intermediate_reg_0[2840]),.o(intermediate_reg_1[1420]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2839]),.i2(intermediate_reg_0[2838]),.o(intermediate_reg_1[1419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2837]),.i2(intermediate_reg_0[2836]),.o(intermediate_reg_1[1418]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2835]),.i2(intermediate_reg_0[2834]),.o(intermediate_reg_1[1417])); 
xor_module xor_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2833]),.i2(intermediate_reg_0[2832]),.o(intermediate_reg_1[1416])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2831]),.i2(intermediate_reg_0[2830]),.o(intermediate_reg_1[1415])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2829]),.i2(intermediate_reg_0[2828]),.o(intermediate_reg_1[1414])); 
xor_module xor_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2827]),.i2(intermediate_reg_0[2826]),.o(intermediate_reg_1[1413])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2825]),.i2(intermediate_reg_0[2824]),.o(intermediate_reg_1[1412])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2823]),.i2(intermediate_reg_0[2822]),.o(intermediate_reg_1[1411]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2821]),.i2(intermediate_reg_0[2820]),.o(intermediate_reg_1[1410]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2819]),.i2(intermediate_reg_0[2818]),.o(intermediate_reg_1[1409]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2817]),.i2(intermediate_reg_0[2816]),.o(intermediate_reg_1[1408])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2815]),.i2(intermediate_reg_0[2814]),.o(intermediate_reg_1[1407])); 
mux_module mux_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2813]),.i2(intermediate_reg_0[2812]),.o(intermediate_reg_1[1406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2811]),.i2(intermediate_reg_0[2810]),.o(intermediate_reg_1[1405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2809]),.i2(intermediate_reg_0[2808]),.o(intermediate_reg_1[1404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2807]),.i2(intermediate_reg_0[2806]),.o(intermediate_reg_1[1403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2805]),.i2(intermediate_reg_0[2804]),.o(intermediate_reg_1[1402]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2803]),.i2(intermediate_reg_0[2802]),.o(intermediate_reg_1[1401])); 
mux_module mux_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2801]),.i2(intermediate_reg_0[2800]),.o(intermediate_reg_1[1400]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2799]),.i2(intermediate_reg_0[2798]),.o(intermediate_reg_1[1399])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2797]),.i2(intermediate_reg_0[2796]),.o(intermediate_reg_1[1398]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2795]),.i2(intermediate_reg_0[2794]),.o(intermediate_reg_1[1397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2793]),.i2(intermediate_reg_0[2792]),.o(intermediate_reg_1[1396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2791]),.i2(intermediate_reg_0[2790]),.o(intermediate_reg_1[1395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2789]),.i2(intermediate_reg_0[2788]),.o(intermediate_reg_1[1394]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2787]),.i2(intermediate_reg_0[2786]),.o(intermediate_reg_1[1393]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2785]),.i2(intermediate_reg_0[2784]),.o(intermediate_reg_1[1392])); 
xor_module xor_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2783]),.i2(intermediate_reg_0[2782]),.o(intermediate_reg_1[1391])); 
xor_module xor_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2781]),.i2(intermediate_reg_0[2780]),.o(intermediate_reg_1[1390])); 
xor_module xor_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2779]),.i2(intermediate_reg_0[2778]),.o(intermediate_reg_1[1389])); 
mux_module mux_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2777]),.i2(intermediate_reg_0[2776]),.o(intermediate_reg_1[1388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2775]),.i2(intermediate_reg_0[2774]),.o(intermediate_reg_1[1387])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2773]),.i2(intermediate_reg_0[2772]),.o(intermediate_reg_1[1386]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2771]),.i2(intermediate_reg_0[2770]),.o(intermediate_reg_1[1385])); 
xor_module xor_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2769]),.i2(intermediate_reg_0[2768]),.o(intermediate_reg_1[1384])); 
mux_module mux_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2767]),.i2(intermediate_reg_0[2766]),.o(intermediate_reg_1[1383]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2765]),.i2(intermediate_reg_0[2764]),.o(intermediate_reg_1[1382])); 
mux_module mux_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2763]),.i2(intermediate_reg_0[2762]),.o(intermediate_reg_1[1381]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2761]),.i2(intermediate_reg_0[2760]),.o(intermediate_reg_1[1380]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2759]),.i2(intermediate_reg_0[2758]),.o(intermediate_reg_1[1379])); 
mux_module mux_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2757]),.i2(intermediate_reg_0[2756]),.o(intermediate_reg_1[1378]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2755]),.i2(intermediate_reg_0[2754]),.o(intermediate_reg_1[1377])); 
xor_module xor_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2753]),.i2(intermediate_reg_0[2752]),.o(intermediate_reg_1[1376])); 
mux_module mux_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2751]),.i2(intermediate_reg_0[2750]),.o(intermediate_reg_1[1375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2749]),.i2(intermediate_reg_0[2748]),.o(intermediate_reg_1[1374]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2747]),.i2(intermediate_reg_0[2746]),.o(intermediate_reg_1[1373])); 
mux_module mux_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2745]),.i2(intermediate_reg_0[2744]),.o(intermediate_reg_1[1372]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2743]),.i2(intermediate_reg_0[2742]),.o(intermediate_reg_1[1371])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2741]),.i2(intermediate_reg_0[2740]),.o(intermediate_reg_1[1370])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2739]),.i2(intermediate_reg_0[2738]),.o(intermediate_reg_1[1369]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2737]),.i2(intermediate_reg_0[2736]),.o(intermediate_reg_1[1368]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2735]),.i2(intermediate_reg_0[2734]),.o(intermediate_reg_1[1367])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2733]),.i2(intermediate_reg_0[2732]),.o(intermediate_reg_1[1366])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2731]),.i2(intermediate_reg_0[2730]),.o(intermediate_reg_1[1365])); 
xor_module xor_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2729]),.i2(intermediate_reg_0[2728]),.o(intermediate_reg_1[1364])); 
mux_module mux_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2727]),.i2(intermediate_reg_0[2726]),.o(intermediate_reg_1[1363]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2725]),.i2(intermediate_reg_0[2724]),.o(intermediate_reg_1[1362]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2723]),.i2(intermediate_reg_0[2722]),.o(intermediate_reg_1[1361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2721]),.i2(intermediate_reg_0[2720]),.o(intermediate_reg_1[1360]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2719]),.i2(intermediate_reg_0[2718]),.o(intermediate_reg_1[1359])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2717]),.i2(intermediate_reg_0[2716]),.o(intermediate_reg_1[1358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2715]),.i2(intermediate_reg_0[2714]),.o(intermediate_reg_1[1357]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2713]),.i2(intermediate_reg_0[2712]),.o(intermediate_reg_1[1356])); 
xor_module xor_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2711]),.i2(intermediate_reg_0[2710]),.o(intermediate_reg_1[1355])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2709]),.i2(intermediate_reg_0[2708]),.o(intermediate_reg_1[1354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2707]),.i2(intermediate_reg_0[2706]),.o(intermediate_reg_1[1353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2705]),.i2(intermediate_reg_0[2704]),.o(intermediate_reg_1[1352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2703]),.i2(intermediate_reg_0[2702]),.o(intermediate_reg_1[1351]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2701]),.i2(intermediate_reg_0[2700]),.o(intermediate_reg_1[1350])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2699]),.i2(intermediate_reg_0[2698]),.o(intermediate_reg_1[1349]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2697]),.i2(intermediate_reg_0[2696]),.o(intermediate_reg_1[1348])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2695]),.i2(intermediate_reg_0[2694]),.o(intermediate_reg_1[1347]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2693]),.i2(intermediate_reg_0[2692]),.o(intermediate_reg_1[1346])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2691]),.i2(intermediate_reg_0[2690]),.o(intermediate_reg_1[1345]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2689]),.i2(intermediate_reg_0[2688]),.o(intermediate_reg_1[1344]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343])); 
mux_module mux_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337])); 
mux_module mux_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332])); 
mux_module mux_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329])); 
mux_module mux_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326])); 
mux_module mux_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320])); 
xor_module xor_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319])); 
mux_module mux_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315])); 
mux_module mux_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311])); 
xor_module xor_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310])); 
mux_module mux_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307])); 
xor_module xor_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302])); 
mux_module mux_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300])); 
mux_module mux_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298])); 
mux_module mux_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295])); 
mux_module mux_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292])); 
mux_module mux_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289])); 
xor_module xor_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286])); 
xor_module xor_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285])); 
xor_module xor_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284])); 
xor_module xor_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283])); 
xor_module xor_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282])); 
xor_module xor_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278])); 
xor_module xor_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277])); 
mux_module mux_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274])); 
xor_module xor_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261])); 
xor_module xor_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260])); 
xor_module xor_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258])); 
xor_module xor_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251])); 
xor_module xor_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246])); 
xor_module xor_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245])); 
xor_module xor_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244])); 
xor_module xor_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241])); 
xor_module xor_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237])); 
xor_module xor_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236])); 
mux_module mux_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232])); 
mux_module mux_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230])); 
mux_module mux_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228])); 
mux_module mux_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
mux_module mux_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224])); 
xor_module xor_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222])); 
xor_module xor_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220])); 
mux_module mux_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218])); 
xor_module xor_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217])); 
xor_module xor_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216])); 
mux_module mux_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211])); 
mux_module mux_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205])); 
xor_module xor_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204])); 
mux_module mux_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202])); 
xor_module xor_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201])); 
xor_module xor_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200])); 
xor_module xor_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199])); 
xor_module xor_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198])); 
mux_module mux_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196])); 
mux_module mux_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194])); 
xor_module xor_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191])); 
xor_module xor_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190])); 
mux_module mux_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183])); 
xor_module xor_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182])); 
mux_module mux_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179])); 
xor_module xor_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178])); 
mux_module mux_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175])); 
mux_module mux_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167])); 
xor_module xor_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166])); 
mux_module mux_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164])); 
xor_module xor_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159])); 
mux_module mux_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156])); 
xor_module xor_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155])); 
mux_module mux_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152])); 
mux_module mux_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145])); 
mux_module mux_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143])); 
xor_module xor_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142])); 
mux_module mux_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137])); 
mux_module mux_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132])); 
mux_module mux_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
mux_module mux_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121])); 
xor_module xor_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120])); 
xor_module xor_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
xor_module xor_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118])); 
xor_module xor_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117])); 
mux_module mux_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115])); 
mux_module mux_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110])); 
mux_module mux_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
xor_module xor_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107])); 
xor_module xor_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106])); 
xor_module xor_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
xor_module xor_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
mux_module mux_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098])); 
mux_module mux_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095])); 
mux_module mux_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
mux_module mux_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
mux_module mux_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082])); 
xor_module xor_module_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081])); 
mux_module mux_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
xor_module xor_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077])); 
mux_module mux_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068])); 
xor_module xor_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
mux_module mux_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064])); 
mux_module mux_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062])); 
mux_module mux_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060])); 
mux_module mux_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058])); 
mux_module mux_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056])); 
mux_module mux_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
mux_module mux_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050])); 
xor_module xor_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049])); 
xor_module xor_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048])); 
xor_module xor_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
xor_module xor_module_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046])); 
mux_module mux_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
xor_module xor_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
xor_module xor_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
mux_module mux_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037])); 
xor_module xor_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036])); 
mux_module mux_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033])); 
mux_module mux_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
mux_module mux_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026])); 
xor_module xor_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
mux_module mux_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021])); 
xor_module xor_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016])); 
xor_module xor_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
xor_module xor_module_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
mux_module mux_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012])); 
xor_module xor_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011])); 
xor_module xor_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010])); 
mux_module mux_module_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
xor_module xor_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
mux_module mux_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
mux_module mux_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
mux_module mux_module_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
mux_module mux_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
mux_module mux_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
xor_module xor_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
mux_module mux_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
xor_module xor_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
mux_module mux_module_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
xor_module xor_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
xor_module xor_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
xor_module xor_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
xor_module xor_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
xor_module xor_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
xor_module xor_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
mux_module mux_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971])); 
mux_module mux_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
mux_module mux_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
xor_module xor_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
xor_module xor_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
mux_module mux_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
xor_module xor_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959])); 
xor_module xor_module_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
mux_module mux_module_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
xor_module xor_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
xor_module xor_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954])); 
mux_module mux_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
mux_module mux_module_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948])); 
xor_module xor_module_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
xor_module xor_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
xor_module xor_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
xor_module xor_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
mux_module mux_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
mux_module mux_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
mux_module mux_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
mux_module mux_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
xor_module xor_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
mux_module mux_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
xor_module xor_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
xor_module xor_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
xor_module xor_module_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
mux_module mux_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
xor_module xor_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
xor_module xor_module_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
mux_module mux_module_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
mux_module mux_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
xor_module xor_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
mux_module mux_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
mux_module mux_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
mux_module mux_module_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
xor_module xor_module_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
xor_module xor_module_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
xor_module xor_module_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
mux_module mux_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
mux_module mux_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
mux_module mux_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
mux_module mux_module_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879])); 
xor_module xor_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
xor_module xor_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
mux_module mux_module_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
mux_module mux_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
mux_module mux_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
xor_module xor_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
xor_module xor_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865])); 
xor_module xor_module_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
mux_module mux_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
xor_module xor_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
xor_module xor_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
xor_module xor_module_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
mux_module mux_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
mux_module mux_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
xor_module xor_module_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
mux_module mux_module_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842])); 
xor_module xor_module_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
mux_module mux_module_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
xor_module xor_module_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
xor_module xor_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
xor_module xor_module_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
mux_module mux_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
mux_module mux_module_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
xor_module xor_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
xor_module xor_module_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
mux_module mux_module_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
xor_module xor_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
mux_module mux_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
xor_module xor_module_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
xor_module xor_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
xor_module xor_module_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
xor_module xor_module_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
mux_module mux_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
xor_module xor_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
mux_module mux_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
xor_module xor_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
xor_module xor_module_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
mux_module mux_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
mux_module mux_module_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
mux_module mux_module_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
xor_module xor_module_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
mux_module mux_module_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
mux_module mux_module_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
xor_module xor_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
xor_module xor_module_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
mux_module mux_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
mux_module mux_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
xor_module xor_module_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
xor_module xor_module_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
mux_module mux_module_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
xor_module xor_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
mux_module mux_module_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
mux_module mux_module_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
xor_module xor_module_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
mux_module mux_module_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
xor_module xor_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
xor_module xor_module_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
xor_module xor_module_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
mux_module mux_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
xor_module xor_module_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
xor_module xor_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
mux_module mux_module_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
mux_module mux_module_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
mux_module mux_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
mux_module mux_module_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
mux_module mux_module_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
mux_module mux_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
xor_module xor_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
mux_module mux_module_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
xor_module xor_module_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
xor_module xor_module_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
xor_module xor_module_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
xor_module xor_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
mux_module mux_module_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
xor_module xor_module_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
mux_module mux_module_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
xor_module xor_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
xor_module xor_module_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
mux_module mux_module_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
xor_module xor_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
xor_module xor_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
xor_module xor_module_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
xor_module xor_module_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
xor_module xor_module_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
xor_module xor_module_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
xor_module xor_module_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
xor_module xor_module_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
xor_module xor_module_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
mux_module mux_module_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
mux_module mux_module_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
xor_module xor_module_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
xor_module xor_module_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
xor_module xor_module_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
xor_module xor_module_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
xor_module xor_module_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
xor_module xor_module_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
mux_module mux_module_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687])); 
mux_module mux_module_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
xor_module xor_module_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
mux_module mux_module_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
xor_module xor_module_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
mux_module mux_module_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
xor_module xor_module_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
mux_module mux_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
mux_module mux_module_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
mux_module mux_module_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
xor_module xor_module_inst_1_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
xor_module xor_module_inst_1_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
mux_module mux_module_inst_1_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
mux_module mux_module_inst_1_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
xor_module xor_module_inst_1_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
mux_module mux_module_inst_1_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
mux_module mux_module_inst_1_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
xor_module xor_module_inst_1_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
mux_module mux_module_inst_1_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
xor_module xor_module_inst_1_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
xor_module xor_module_inst_1_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
xor_module xor_module_inst_1_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
xor_module xor_module_inst_1_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
xor_module xor_module_inst_1_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642])); 
mux_module mux_module_inst_1_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
xor_module xor_module_inst_1_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
xor_module xor_module_inst_1_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
mux_module mux_module_inst_1_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
xor_module xor_module_inst_1_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
xor_module xor_module_inst_1_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
mux_module mux_module_inst_1_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
xor_module xor_module_inst_1_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
xor_module xor_module_inst_1_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
xor_module xor_module_inst_1_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
xor_module xor_module_inst_1_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
mux_module mux_module_inst_1_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
mux_module mux_module_inst_1_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
xor_module xor_module_inst_1_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
mux_module mux_module_inst_1_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
xor_module xor_module_inst_1_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
xor_module xor_module_inst_1_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
xor_module xor_module_inst_1_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
mux_module mux_module_inst_1_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
xor_module xor_module_inst_1_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
xor_module xor_module_inst_1_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
xor_module xor_module_inst_1_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
mux_module mux_module_inst_1_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
xor_module xor_module_inst_1_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
xor_module xor_module_inst_1_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
mux_module mux_module_inst_1_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
xor_module xor_module_inst_1_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
mux_module mux_module_inst_1_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
mux_module mux_module_inst_1_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
mux_module mux_module_inst_1_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
mux_module mux_module_inst_1_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
mux_module mux_module_inst_1_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
xor_module xor_module_inst_1_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
xor_module xor_module_inst_1_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
mux_module mux_module_inst_1_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
xor_module xor_module_inst_1_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
mux_module mux_module_inst_1_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
xor_module xor_module_inst_1_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
xor_module xor_module_inst_1_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
mux_module mux_module_inst_1_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
mux_module mux_module_inst_1_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
xor_module xor_module_inst_1_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
xor_module xor_module_inst_1_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
xor_module xor_module_inst_1_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
mux_module mux_module_inst_1_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
mux_module mux_module_inst_1_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
mux_module mux_module_inst_1_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
xor_module xor_module_inst_1_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
mux_module mux_module_inst_1_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
xor_module xor_module_inst_1_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
xor_module xor_module_inst_1_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
xor_module xor_module_inst_1_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
mux_module mux_module_inst_1_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
xor_module xor_module_inst_1_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
xor_module xor_module_inst_1_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
mux_module mux_module_inst_1_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
xor_module xor_module_inst_1_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
mux_module mux_module_inst_1_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
mux_module mux_module_inst_1_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
mux_module mux_module_inst_1_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
xor_module xor_module_inst_1_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
mux_module mux_module_inst_1_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
xor_module xor_module_inst_1_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
mux_module mux_module_inst_1_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
mux_module mux_module_inst_1_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
xor_module xor_module_inst_1_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
xor_module xor_module_inst_1_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
xor_module xor_module_inst_1_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
mux_module mux_module_inst_1_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
mux_module mux_module_inst_1_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
mux_module mux_module_inst_1_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
xor_module xor_module_inst_1_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
xor_module xor_module_inst_1_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
mux_module mux_module_inst_1_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
mux_module mux_module_inst_1_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
mux_module mux_module_inst_1_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
mux_module mux_module_inst_1_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
mux_module mux_module_inst_1_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
xor_module xor_module_inst_1_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
xor_module xor_module_inst_1_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
xor_module xor_module_inst_1_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
mux_module mux_module_inst_1_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
xor_module xor_module_inst_1_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
mux_module mux_module_inst_1_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
xor_module xor_module_inst_1_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
mux_module mux_module_inst_1_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
mux_module mux_module_inst_1_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
xor_module xor_module_inst_1_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
mux_module mux_module_inst_1_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
mux_module mux_module_inst_1_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
xor_module xor_module_inst_1_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
mux_module mux_module_inst_1_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
mux_module mux_module_inst_1_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
mux_module mux_module_inst_1_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
xor_module xor_module_inst_1_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
mux_module mux_module_inst_1_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
mux_module mux_module_inst_1_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
xor_module xor_module_inst_1_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
xor_module xor_module_inst_1_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
xor_module xor_module_inst_1_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
mux_module mux_module_inst_1_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
xor_module xor_module_inst_1_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
mux_module mux_module_inst_1_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
xor_module xor_module_inst_1_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
xor_module xor_module_inst_1_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
xor_module xor_module_inst_1_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
xor_module xor_module_inst_1_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
xor_module xor_module_inst_1_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
mux_module mux_module_inst_1_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
mux_module mux_module_inst_1_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
xor_module xor_module_inst_1_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
xor_module xor_module_inst_1_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
mux_module mux_module_inst_1_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
xor_module xor_module_inst_1_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
mux_module mux_module_inst_1_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
xor_module xor_module_inst_1_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
mux_module mux_module_inst_1_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
xor_module xor_module_inst_1_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
mux_module mux_module_inst_1_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
mux_module mux_module_inst_1_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
xor_module xor_module_inst_1_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
mux_module mux_module_inst_1_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
mux_module mux_module_inst_1_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
xor_module xor_module_inst_1_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
xor_module xor_module_inst_1_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
mux_module mux_module_inst_1_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
mux_module mux_module_inst_1_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
xor_module xor_module_inst_1_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
mux_module mux_module_inst_1_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
xor_module xor_module_inst_1_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
xor_module xor_module_inst_1_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
mux_module mux_module_inst_1_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
xor_module xor_module_inst_1_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
xor_module xor_module_inst_1_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
xor_module xor_module_inst_1_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
mux_module mux_module_inst_1_1649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
xor_module xor_module_inst_1_1653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
mux_module mux_module_inst_1_1654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
xor_module xor_module_inst_1_1657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
xor_module xor_module_inst_1_1658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
mux_module mux_module_inst_1_1659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
mux_module mux_module_inst_1_1661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
xor_module xor_module_inst_1_1664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
mux_module mux_module_inst_1_1665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
mux_module mux_module_inst_1_1668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
xor_module xor_module_inst_1_1670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
mux_module mux_module_inst_1_1671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
xor_module xor_module_inst_1_1673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
mux_module mux_module_inst_1_1674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
mux_module mux_module_inst_1_1676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
mux_module mux_module_inst_1_1678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
xor_module xor_module_inst_1_1681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_1682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
mux_module mux_module_inst_1_1683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
mux_module mux_module_inst_1_1685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_1687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
xor_module xor_module_inst_1_1688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
mux_module mux_module_inst_1_1689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
xor_module xor_module_inst_1_1692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
xor_module xor_module_inst_1_1693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
xor_module xor_module_inst_1_1694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
xor_module xor_module_inst_1_1695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
xor_module xor_module_inst_1_1696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_1697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
mux_module mux_module_inst_1_1700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
xor_module xor_module_inst_1_1702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
mux_module mux_module_inst_1_1703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
xor_module xor_module_inst_1_1708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
xor_module xor_module_inst_1_1709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
xor_module xor_module_inst_1_1710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
mux_module mux_module_inst_1_1711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
mux_module mux_module_inst_1_1713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
xor_module xor_module_inst_1_1721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
mux_module mux_module_inst_1_1722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
xor_module xor_module_inst_1_1725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
xor_module xor_module_inst_1_1726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
xor_module xor_module_inst_1_1727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
mux_module mux_module_inst_1_1728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
mux_module mux_module_inst_1_1730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
xor_module xor_module_inst_1_1732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
xor_module xor_module_inst_1_1733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
mux_module mux_module_inst_1_1734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
xor_module xor_module_inst_1_1737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
mux_module mux_module_inst_1_1738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
mux_module mux_module_inst_1_1740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
xor_module xor_module_inst_1_1744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
mux_module mux_module_inst_1_1745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
xor_module xor_module_inst_1_1750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
xor_module xor_module_inst_1_1751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
xor_module xor_module_inst_1_1752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
mux_module mux_module_inst_1_1753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
mux_module mux_module_inst_1_1755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
xor_module xor_module_inst_1_1759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_1760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
mux_module mux_module_inst_1_1761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
mux_module mux_module_inst_1_1765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
mux_module mux_module_inst_1_1768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
mux_module mux_module_inst_1_1770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
xor_module xor_module_inst_1_1772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_1773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
xor_module xor_module_inst_1_1774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
mux_module mux_module_inst_1_1775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
mux_module mux_module_inst_1_1777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
mux_module mux_module_inst_1_1779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
mux_module mux_module_inst_1_1781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
xor_module xor_module_inst_1_1786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
xor_module xor_module_inst_1_1787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
mux_module mux_module_inst_1_1788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_1790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_1791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
xor_module xor_module_inst_1_1792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
xor_module xor_module_inst_1_1793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
xor_module xor_module_inst_1_1794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
xor_module xor_module_inst_1_1795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
xor_module xor_module_inst_1_1796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
mux_module mux_module_inst_1_1797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
xor_module xor_module_inst_1_1800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
xor_module xor_module_inst_1_1801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
xor_module xor_module_inst_1_1802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
mux_module mux_module_inst_1_1803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
mux_module mux_module_inst_1_1807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_1810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
xor_module xor_module_inst_1_1813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
mux_module mux_module_inst_1_1814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
mux_module mux_module_inst_1_1817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
mux_module mux_module_inst_1_1821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
mux_module mux_module_inst_1_1824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
mux_module mux_module_inst_1_1827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
xor_module xor_module_inst_1_1830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_1831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
xor_module xor_module_inst_1_1832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
mux_module mux_module_inst_1_1833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
xor_module xor_module_inst_1_1835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
xor_module xor_module_inst_1_1836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
mux_module mux_module_inst_1_1837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
mux_module mux_module_inst_1_1840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
xor_module xor_module_inst_1_1842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
xor_module xor_module_inst_1_1843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
xor_module xor_module_inst_1_1844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
xor_module xor_module_inst_1_1845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
mux_module mux_module_inst_1_1846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
xor_module xor_module_inst_1_1848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
xor_module xor_module_inst_1_1849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_1850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
mux_module mux_module_inst_1_1851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_1853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
xor_module xor_module_inst_1_1854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
mux_module mux_module_inst_1_1855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
xor_module xor_module_inst_1_1857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
xor_module xor_module_inst_1_1858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
mux_module mux_module_inst_1_1859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
mux_module mux_module_inst_1_1862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_1864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
xor_module xor_module_inst_1_1865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
mux_module mux_module_inst_1_1866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
xor_module xor_module_inst_1_1868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
mux_module mux_module_inst_1_1869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
mux_module mux_module_inst_1_1872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
xor_module xor_module_inst_1_1874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
mux_module mux_module_inst_1_1875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
mux_module mux_module_inst_1_1879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
mux_module mux_module_inst_1_1881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
xor_module xor_module_inst_1_1884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
mux_module mux_module_inst_1_1885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
xor_module xor_module_inst_1_1887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
xor_module xor_module_inst_1_1888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
mux_module mux_module_inst_1_1889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_1893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
mux_module mux_module_inst_1_1894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
mux_module mux_module_inst_1_1897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
mux_module mux_module_inst_1_1900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_1903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
xor_module xor_module_inst_1_1904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
mux_module mux_module_inst_1_1905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
mux_module mux_module_inst_1_1907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
mux_module mux_module_inst_1_1911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_1914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
xor_module xor_module_inst_1_1918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
xor_module xor_module_inst_1_1919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
mux_module mux_module_inst_1_1920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
mux_module mux_module_inst_1_1922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
mux_module mux_module_inst_1_1925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
xor_module xor_module_inst_1_1927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
xor_module xor_module_inst_1_1928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
xor_module xor_module_inst_1_1929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
mux_module mux_module_inst_1_1930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
mux_module mux_module_inst_1_1933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
xor_module xor_module_inst_1_1935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
mux_module mux_module_inst_1_1936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_1938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
xor_module xor_module_inst_1_1940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_1941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_1942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
mux_module mux_module_inst_1_1944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
xor_module xor_module_inst_1_1946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
mux_module mux_module_inst_1_1947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
xor_module xor_module_inst_1_1950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
xor_module xor_module_inst_1_1951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
mux_module mux_module_inst_1_1952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
xor_module xor_module_inst_1_1954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
mux_module mux_module_inst_1_1955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
mux_module mux_module_inst_1_1957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
mux_module mux_module_inst_1_1959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
mux_module mux_module_inst_1_1961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
xor_module xor_module_inst_1_1966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_1967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
mux_module mux_module_inst_1_1972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_1974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_1975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
mux_module mux_module_inst_1_1976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
mux_module mux_module_inst_1_1978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
mux_module mux_module_inst_1_1980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
mux_module mux_module_inst_1_1982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_1985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
xor_module xor_module_inst_1_1986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
xor_module xor_module_inst_1_1987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
xor_module xor_module_inst_1_1988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
xor_module xor_module_inst_1_1989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
xor_module xor_module_inst_1_1990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
mux_module mux_module_inst_1_1991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
xor_module xor_module_inst_1_1997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
xor_module xor_module_inst_1_1998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
xor_module xor_module_inst_1_1999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
mux_module mux_module_inst_1_2000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_2004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
mux_module mux_module_inst_1_2005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
reg [1003:0]intermediate_reg_2; 
 
xor_module xor_module_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2007]),.i2(intermediate_reg_1[2006]),.o(intermediate_reg_2[1003])); 
xor_module xor_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2005]),.i2(intermediate_reg_1[2004]),.o(intermediate_reg_2[1002])); 
mux_module mux_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2003]),.i2(intermediate_reg_1[2002]),.o(intermediate_reg_2[1001]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2001]),.i2(intermediate_reg_1[2000]),.o(intermediate_reg_2[1000]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1999]),.i2(intermediate_reg_1[1998]),.o(intermediate_reg_2[999])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1997]),.i2(intermediate_reg_1[1996]),.o(intermediate_reg_2[998]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1995]),.i2(intermediate_reg_1[1994]),.o(intermediate_reg_2[997]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1993]),.i2(intermediate_reg_1[1992]),.o(intermediate_reg_2[996])); 
mux_module mux_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1991]),.i2(intermediate_reg_1[1990]),.o(intermediate_reg_2[995]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1989]),.i2(intermediate_reg_1[1988]),.o(intermediate_reg_2[994])); 
mux_module mux_module_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1987]),.i2(intermediate_reg_1[1986]),.o(intermediate_reg_2[993]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1985]),.i2(intermediate_reg_1[1984]),.o(intermediate_reg_2[992]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1983]),.i2(intermediate_reg_1[1982]),.o(intermediate_reg_2[991]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1981]),.i2(intermediate_reg_1[1980]),.o(intermediate_reg_2[990]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1979]),.i2(intermediate_reg_1[1978]),.o(intermediate_reg_2[989])); 
xor_module xor_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1977]),.i2(intermediate_reg_1[1976]),.o(intermediate_reg_2[988])); 
xor_module xor_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1975]),.i2(intermediate_reg_1[1974]),.o(intermediate_reg_2[987])); 
xor_module xor_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1973]),.i2(intermediate_reg_1[1972]),.o(intermediate_reg_2[986])); 
mux_module mux_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1971]),.i2(intermediate_reg_1[1970]),.o(intermediate_reg_2[985]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1969]),.i2(intermediate_reg_1[1968]),.o(intermediate_reg_2[984])); 
xor_module xor_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1967]),.i2(intermediate_reg_1[1966]),.o(intermediate_reg_2[983])); 
xor_module xor_module_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1965]),.i2(intermediate_reg_1[1964]),.o(intermediate_reg_2[982])); 
xor_module xor_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1963]),.i2(intermediate_reg_1[1962]),.o(intermediate_reg_2[981])); 
mux_module mux_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1961]),.i2(intermediate_reg_1[1960]),.o(intermediate_reg_2[980]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1959]),.i2(intermediate_reg_1[1958]),.o(intermediate_reg_2[979])); 
mux_module mux_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1957]),.i2(intermediate_reg_1[1956]),.o(intermediate_reg_2[978]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1955]),.i2(intermediate_reg_1[1954]),.o(intermediate_reg_2[977])); 
xor_module xor_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1953]),.i2(intermediate_reg_1[1952]),.o(intermediate_reg_2[976])); 
mux_module mux_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1951]),.i2(intermediate_reg_1[1950]),.o(intermediate_reg_2[975]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1949]),.i2(intermediate_reg_1[1948]),.o(intermediate_reg_2[974])); 
xor_module xor_module_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1947]),.i2(intermediate_reg_1[1946]),.o(intermediate_reg_2[973])); 
mux_module mux_module_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1945]),.i2(intermediate_reg_1[1944]),.o(intermediate_reg_2[972]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1943]),.i2(intermediate_reg_1[1942]),.o(intermediate_reg_2[971])); 
xor_module xor_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1941]),.i2(intermediate_reg_1[1940]),.o(intermediate_reg_2[970])); 
xor_module xor_module_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1939]),.i2(intermediate_reg_1[1938]),.o(intermediate_reg_2[969])); 
xor_module xor_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1937]),.i2(intermediate_reg_1[1936]),.o(intermediate_reg_2[968])); 
xor_module xor_module_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1935]),.i2(intermediate_reg_1[1934]),.o(intermediate_reg_2[967])); 
mux_module mux_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1933]),.i2(intermediate_reg_1[1932]),.o(intermediate_reg_2[966]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1931]),.i2(intermediate_reg_1[1930]),.o(intermediate_reg_2[965]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1929]),.i2(intermediate_reg_1[1928]),.o(intermediate_reg_2[964])); 
mux_module mux_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1927]),.i2(intermediate_reg_1[1926]),.o(intermediate_reg_2[963]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1925]),.i2(intermediate_reg_1[1924]),.o(intermediate_reg_2[962]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1923]),.i2(intermediate_reg_1[1922]),.o(intermediate_reg_2[961])); 
xor_module xor_module_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1921]),.i2(intermediate_reg_1[1920]),.o(intermediate_reg_2[960])); 
xor_module xor_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1919]),.i2(intermediate_reg_1[1918]),.o(intermediate_reg_2[959])); 
mux_module mux_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1917]),.i2(intermediate_reg_1[1916]),.o(intermediate_reg_2[958]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1915]),.i2(intermediate_reg_1[1914]),.o(intermediate_reg_2[957])); 
mux_module mux_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1913]),.i2(intermediate_reg_1[1912]),.o(intermediate_reg_2[956]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1911]),.i2(intermediate_reg_1[1910]),.o(intermediate_reg_2[955])); 
xor_module xor_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1909]),.i2(intermediate_reg_1[1908]),.o(intermediate_reg_2[954])); 
xor_module xor_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1907]),.i2(intermediate_reg_1[1906]),.o(intermediate_reg_2[953])); 
xor_module xor_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1905]),.i2(intermediate_reg_1[1904]),.o(intermediate_reg_2[952])); 
mux_module mux_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1903]),.i2(intermediate_reg_1[1902]),.o(intermediate_reg_2[951]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1901]),.i2(intermediate_reg_1[1900]),.o(intermediate_reg_2[950])); 
xor_module xor_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1899]),.i2(intermediate_reg_1[1898]),.o(intermediate_reg_2[949])); 
xor_module xor_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1897]),.i2(intermediate_reg_1[1896]),.o(intermediate_reg_2[948])); 
mux_module mux_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1895]),.i2(intermediate_reg_1[1894]),.o(intermediate_reg_2[947]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1893]),.i2(intermediate_reg_1[1892]),.o(intermediate_reg_2[946])); 
mux_module mux_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1891]),.i2(intermediate_reg_1[1890]),.o(intermediate_reg_2[945]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1889]),.i2(intermediate_reg_1[1888]),.o(intermediate_reg_2[944]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1887]),.i2(intermediate_reg_1[1886]),.o(intermediate_reg_2[943]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1885]),.i2(intermediate_reg_1[1884]),.o(intermediate_reg_2[942])); 
mux_module mux_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1883]),.i2(intermediate_reg_1[1882]),.o(intermediate_reg_2[941]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1881]),.i2(intermediate_reg_1[1880]),.o(intermediate_reg_2[940]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1879]),.i2(intermediate_reg_1[1878]),.o(intermediate_reg_2[939])); 
mux_module mux_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1877]),.i2(intermediate_reg_1[1876]),.o(intermediate_reg_2[938]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1875]),.i2(intermediate_reg_1[1874]),.o(intermediate_reg_2[937])); 
mux_module mux_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1873]),.i2(intermediate_reg_1[1872]),.o(intermediate_reg_2[936]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1871]),.i2(intermediate_reg_1[1870]),.o(intermediate_reg_2[935])); 
xor_module xor_module_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1869]),.i2(intermediate_reg_1[1868]),.o(intermediate_reg_2[934])); 
xor_module xor_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1867]),.i2(intermediate_reg_1[1866]),.o(intermediate_reg_2[933])); 
mux_module mux_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1865]),.i2(intermediate_reg_1[1864]),.o(intermediate_reg_2[932]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1863]),.i2(intermediate_reg_1[1862]),.o(intermediate_reg_2[931]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1861]),.i2(intermediate_reg_1[1860]),.o(intermediate_reg_2[930]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1859]),.i2(intermediate_reg_1[1858]),.o(intermediate_reg_2[929])); 
mux_module mux_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1857]),.i2(intermediate_reg_1[1856]),.o(intermediate_reg_2[928]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1855]),.i2(intermediate_reg_1[1854]),.o(intermediate_reg_2[927]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1853]),.i2(intermediate_reg_1[1852]),.o(intermediate_reg_2[926]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1851]),.i2(intermediate_reg_1[1850]),.o(intermediate_reg_2[925])); 
mux_module mux_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1849]),.i2(intermediate_reg_1[1848]),.o(intermediate_reg_2[924]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1847]),.i2(intermediate_reg_1[1846]),.o(intermediate_reg_2[923])); 
xor_module xor_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1845]),.i2(intermediate_reg_1[1844]),.o(intermediate_reg_2[922])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1843]),.i2(intermediate_reg_1[1842]),.o(intermediate_reg_2[921]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1841]),.i2(intermediate_reg_1[1840]),.o(intermediate_reg_2[920])); 
xor_module xor_module_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1839]),.i2(intermediate_reg_1[1838]),.o(intermediate_reg_2[919])); 
xor_module xor_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1837]),.i2(intermediate_reg_1[1836]),.o(intermediate_reg_2[918])); 
mux_module mux_module_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1835]),.i2(intermediate_reg_1[1834]),.o(intermediate_reg_2[917]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1833]),.i2(intermediate_reg_1[1832]),.o(intermediate_reg_2[916]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1831]),.i2(intermediate_reg_1[1830]),.o(intermediate_reg_2[915])); 
xor_module xor_module_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1829]),.i2(intermediate_reg_1[1828]),.o(intermediate_reg_2[914])); 
xor_module xor_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1827]),.i2(intermediate_reg_1[1826]),.o(intermediate_reg_2[913])); 
xor_module xor_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1825]),.i2(intermediate_reg_1[1824]),.o(intermediate_reg_2[912])); 
xor_module xor_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1823]),.i2(intermediate_reg_1[1822]),.o(intermediate_reg_2[911])); 
mux_module mux_module_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1821]),.i2(intermediate_reg_1[1820]),.o(intermediate_reg_2[910]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1819]),.i2(intermediate_reg_1[1818]),.o(intermediate_reg_2[909]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1817]),.i2(intermediate_reg_1[1816]),.o(intermediate_reg_2[908])); 
xor_module xor_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1815]),.i2(intermediate_reg_1[1814]),.o(intermediate_reg_2[907])); 
xor_module xor_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1813]),.i2(intermediate_reg_1[1812]),.o(intermediate_reg_2[906])); 
mux_module mux_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1811]),.i2(intermediate_reg_1[1810]),.o(intermediate_reg_2[905]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1809]),.i2(intermediate_reg_1[1808]),.o(intermediate_reg_2[904]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1807]),.i2(intermediate_reg_1[1806]),.o(intermediate_reg_2[903]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1805]),.i2(intermediate_reg_1[1804]),.o(intermediate_reg_2[902]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1803]),.i2(intermediate_reg_1[1802]),.o(intermediate_reg_2[901])); 
xor_module xor_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1801]),.i2(intermediate_reg_1[1800]),.o(intermediate_reg_2[900])); 
mux_module mux_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1799]),.i2(intermediate_reg_1[1798]),.o(intermediate_reg_2[899]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1797]),.i2(intermediate_reg_1[1796]),.o(intermediate_reg_2[898])); 
xor_module xor_module_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1795]),.i2(intermediate_reg_1[1794]),.o(intermediate_reg_2[897])); 
xor_module xor_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1793]),.i2(intermediate_reg_1[1792]),.o(intermediate_reg_2[896])); 
mux_module mux_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1791]),.i2(intermediate_reg_1[1790]),.o(intermediate_reg_2[895]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1789]),.i2(intermediate_reg_1[1788]),.o(intermediate_reg_2[894]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1787]),.i2(intermediate_reg_1[1786]),.o(intermediate_reg_2[893]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1785]),.i2(intermediate_reg_1[1784]),.o(intermediate_reg_2[892]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1783]),.i2(intermediate_reg_1[1782]),.o(intermediate_reg_2[891])); 
xor_module xor_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1781]),.i2(intermediate_reg_1[1780]),.o(intermediate_reg_2[890])); 
xor_module xor_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1779]),.i2(intermediate_reg_1[1778]),.o(intermediate_reg_2[889])); 
mux_module mux_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1777]),.i2(intermediate_reg_1[1776]),.o(intermediate_reg_2[888]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1775]),.i2(intermediate_reg_1[1774]),.o(intermediate_reg_2[887])); 
xor_module xor_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1773]),.i2(intermediate_reg_1[1772]),.o(intermediate_reg_2[886])); 
xor_module xor_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1771]),.i2(intermediate_reg_1[1770]),.o(intermediate_reg_2[885])); 
xor_module xor_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1769]),.i2(intermediate_reg_1[1768]),.o(intermediate_reg_2[884])); 
mux_module mux_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1767]),.i2(intermediate_reg_1[1766]),.o(intermediate_reg_2[883]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1765]),.i2(intermediate_reg_1[1764]),.o(intermediate_reg_2[882])); 
xor_module xor_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1763]),.i2(intermediate_reg_1[1762]),.o(intermediate_reg_2[881])); 
mux_module mux_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1761]),.i2(intermediate_reg_1[1760]),.o(intermediate_reg_2[880]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1759]),.i2(intermediate_reg_1[1758]),.o(intermediate_reg_2[879])); 
mux_module mux_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1757]),.i2(intermediate_reg_1[1756]),.o(intermediate_reg_2[878]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1755]),.i2(intermediate_reg_1[1754]),.o(intermediate_reg_2[877]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1753]),.i2(intermediate_reg_1[1752]),.o(intermediate_reg_2[876]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1751]),.i2(intermediate_reg_1[1750]),.o(intermediate_reg_2[875])); 
xor_module xor_module_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1749]),.i2(intermediate_reg_1[1748]),.o(intermediate_reg_2[874])); 
mux_module mux_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1747]),.i2(intermediate_reg_1[1746]),.o(intermediate_reg_2[873]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1745]),.i2(intermediate_reg_1[1744]),.o(intermediate_reg_2[872])); 
xor_module xor_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1743]),.i2(intermediate_reg_1[1742]),.o(intermediate_reg_2[871])); 
xor_module xor_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1741]),.i2(intermediate_reg_1[1740]),.o(intermediate_reg_2[870])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1739]),.i2(intermediate_reg_1[1738]),.o(intermediate_reg_2[869]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1737]),.i2(intermediate_reg_1[1736]),.o(intermediate_reg_2[868]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1735]),.i2(intermediate_reg_1[1734]),.o(intermediate_reg_2[867]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1733]),.i2(intermediate_reg_1[1732]),.o(intermediate_reg_2[866])); 
mux_module mux_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1731]),.i2(intermediate_reg_1[1730]),.o(intermediate_reg_2[865]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1729]),.i2(intermediate_reg_1[1728]),.o(intermediate_reg_2[864])); 
xor_module xor_module_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1727]),.i2(intermediate_reg_1[1726]),.o(intermediate_reg_2[863])); 
mux_module mux_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1725]),.i2(intermediate_reg_1[1724]),.o(intermediate_reg_2[862]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1723]),.i2(intermediate_reg_1[1722]),.o(intermediate_reg_2[861])); 
mux_module mux_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1721]),.i2(intermediate_reg_1[1720]),.o(intermediate_reg_2[860]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1719]),.i2(intermediate_reg_1[1718]),.o(intermediate_reg_2[859])); 
mux_module mux_module_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1717]),.i2(intermediate_reg_1[1716]),.o(intermediate_reg_2[858]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1715]),.i2(intermediate_reg_1[1714]),.o(intermediate_reg_2[857])); 
mux_module mux_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1713]),.i2(intermediate_reg_1[1712]),.o(intermediate_reg_2[856]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1711]),.i2(intermediate_reg_1[1710]),.o(intermediate_reg_2[855]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1709]),.i2(intermediate_reg_1[1708]),.o(intermediate_reg_2[854]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1707]),.i2(intermediate_reg_1[1706]),.o(intermediate_reg_2[853]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1705]),.i2(intermediate_reg_1[1704]),.o(intermediate_reg_2[852]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1703]),.i2(intermediate_reg_1[1702]),.o(intermediate_reg_2[851])); 
mux_module mux_module_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1701]),.i2(intermediate_reg_1[1700]),.o(intermediate_reg_2[850]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1699]),.i2(intermediate_reg_1[1698]),.o(intermediate_reg_2[849])); 
mux_module mux_module_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1697]),.i2(intermediate_reg_1[1696]),.o(intermediate_reg_2[848]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1695]),.i2(intermediate_reg_1[1694]),.o(intermediate_reg_2[847]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1693]),.i2(intermediate_reg_1[1692]),.o(intermediate_reg_2[846]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1691]),.i2(intermediate_reg_1[1690]),.o(intermediate_reg_2[845]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1689]),.i2(intermediate_reg_1[1688]),.o(intermediate_reg_2[844])); 
xor_module xor_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1687]),.i2(intermediate_reg_1[1686]),.o(intermediate_reg_2[843])); 
xor_module xor_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1685]),.i2(intermediate_reg_1[1684]),.o(intermediate_reg_2[842])); 
xor_module xor_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1683]),.i2(intermediate_reg_1[1682]),.o(intermediate_reg_2[841])); 
xor_module xor_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1681]),.i2(intermediate_reg_1[1680]),.o(intermediate_reg_2[840])); 
mux_module mux_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1679]),.i2(intermediate_reg_1[1678]),.o(intermediate_reg_2[839]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1677]),.i2(intermediate_reg_1[1676]),.o(intermediate_reg_2[838])); 
mux_module mux_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1675]),.i2(intermediate_reg_1[1674]),.o(intermediate_reg_2[837]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1673]),.i2(intermediate_reg_1[1672]),.o(intermediate_reg_2[836])); 
mux_module mux_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1671]),.i2(intermediate_reg_1[1670]),.o(intermediate_reg_2[835]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1669]),.i2(intermediate_reg_1[1668]),.o(intermediate_reg_2[834]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1667]),.i2(intermediate_reg_1[1666]),.o(intermediate_reg_2[833])); 
xor_module xor_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1665]),.i2(intermediate_reg_1[1664]),.o(intermediate_reg_2[832])); 
mux_module mux_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1663]),.i2(intermediate_reg_1[1662]),.o(intermediate_reg_2[831]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1661]),.i2(intermediate_reg_1[1660]),.o(intermediate_reg_2[830])); 
mux_module mux_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1659]),.i2(intermediate_reg_1[1658]),.o(intermediate_reg_2[829]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1657]),.i2(intermediate_reg_1[1656]),.o(intermediate_reg_2[828]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1655]),.i2(intermediate_reg_1[1654]),.o(intermediate_reg_2[827]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1653]),.i2(intermediate_reg_1[1652]),.o(intermediate_reg_2[826])); 
xor_module xor_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1651]),.i2(intermediate_reg_1[1650]),.o(intermediate_reg_2[825])); 
mux_module mux_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1649]),.i2(intermediate_reg_1[1648]),.o(intermediate_reg_2[824]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1647]),.i2(intermediate_reg_1[1646]),.o(intermediate_reg_2[823]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1645]),.i2(intermediate_reg_1[1644]),.o(intermediate_reg_2[822])); 
mux_module mux_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1643]),.i2(intermediate_reg_1[1642]),.o(intermediate_reg_2[821]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1641]),.i2(intermediate_reg_1[1640]),.o(intermediate_reg_2[820])); 
xor_module xor_module_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1639]),.i2(intermediate_reg_1[1638]),.o(intermediate_reg_2[819])); 
mux_module mux_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1637]),.i2(intermediate_reg_1[1636]),.o(intermediate_reg_2[818]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1635]),.i2(intermediate_reg_1[1634]),.o(intermediate_reg_2[817])); 
mux_module mux_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1633]),.i2(intermediate_reg_1[1632]),.o(intermediate_reg_2[816]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1631]),.i2(intermediate_reg_1[1630]),.o(intermediate_reg_2[815]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1629]),.i2(intermediate_reg_1[1628]),.o(intermediate_reg_2[814])); 
xor_module xor_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1627]),.i2(intermediate_reg_1[1626]),.o(intermediate_reg_2[813])); 
mux_module mux_module_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1625]),.i2(intermediate_reg_1[1624]),.o(intermediate_reg_2[812]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1623]),.i2(intermediate_reg_1[1622]),.o(intermediate_reg_2[811])); 
mux_module mux_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1621]),.i2(intermediate_reg_1[1620]),.o(intermediate_reg_2[810]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1619]),.i2(intermediate_reg_1[1618]),.o(intermediate_reg_2[809]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1617]),.i2(intermediate_reg_1[1616]),.o(intermediate_reg_2[808]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1615]),.i2(intermediate_reg_1[1614]),.o(intermediate_reg_2[807]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1613]),.i2(intermediate_reg_1[1612]),.o(intermediate_reg_2[806]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1611]),.i2(intermediate_reg_1[1610]),.o(intermediate_reg_2[805])); 
xor_module xor_module_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1609]),.i2(intermediate_reg_1[1608]),.o(intermediate_reg_2[804])); 
mux_module mux_module_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1607]),.i2(intermediate_reg_1[1606]),.o(intermediate_reg_2[803]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1605]),.i2(intermediate_reg_1[1604]),.o(intermediate_reg_2[802]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1603]),.i2(intermediate_reg_1[1602]),.o(intermediate_reg_2[801]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1601]),.i2(intermediate_reg_1[1600]),.o(intermediate_reg_2[800])); 
mux_module mux_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1599]),.i2(intermediate_reg_1[1598]),.o(intermediate_reg_2[799]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1597]),.i2(intermediate_reg_1[1596]),.o(intermediate_reg_2[798]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1595]),.i2(intermediate_reg_1[1594]),.o(intermediate_reg_2[797]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1593]),.i2(intermediate_reg_1[1592]),.o(intermediate_reg_2[796])); 
xor_module xor_module_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1591]),.i2(intermediate_reg_1[1590]),.o(intermediate_reg_2[795])); 
mux_module mux_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1589]),.i2(intermediate_reg_1[1588]),.o(intermediate_reg_2[794]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1587]),.i2(intermediate_reg_1[1586]),.o(intermediate_reg_2[793])); 
xor_module xor_module_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1585]),.i2(intermediate_reg_1[1584]),.o(intermediate_reg_2[792])); 
mux_module mux_module_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1583]),.i2(intermediate_reg_1[1582]),.o(intermediate_reg_2[791]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1581]),.i2(intermediate_reg_1[1580]),.o(intermediate_reg_2[790])); 
xor_module xor_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1579]),.i2(intermediate_reg_1[1578]),.o(intermediate_reg_2[789])); 
mux_module mux_module_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1577]),.i2(intermediate_reg_1[1576]),.o(intermediate_reg_2[788]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1575]),.i2(intermediate_reg_1[1574]),.o(intermediate_reg_2[787]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1573]),.i2(intermediate_reg_1[1572]),.o(intermediate_reg_2[786])); 
xor_module xor_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1571]),.i2(intermediate_reg_1[1570]),.o(intermediate_reg_2[785])); 
mux_module mux_module_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1569]),.i2(intermediate_reg_1[1568]),.o(intermediate_reg_2[784]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1567]),.i2(intermediate_reg_1[1566]),.o(intermediate_reg_2[783])); 
mux_module mux_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1565]),.i2(intermediate_reg_1[1564]),.o(intermediate_reg_2[782]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1563]),.i2(intermediate_reg_1[1562]),.o(intermediate_reg_2[781])); 
mux_module mux_module_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1561]),.i2(intermediate_reg_1[1560]),.o(intermediate_reg_2[780]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1559]),.i2(intermediate_reg_1[1558]),.o(intermediate_reg_2[779]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1557]),.i2(intermediate_reg_1[1556]),.o(intermediate_reg_2[778]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1555]),.i2(intermediate_reg_1[1554]),.o(intermediate_reg_2[777]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1553]),.i2(intermediate_reg_1[1552]),.o(intermediate_reg_2[776])); 
xor_module xor_module_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1551]),.i2(intermediate_reg_1[1550]),.o(intermediate_reg_2[775])); 
xor_module xor_module_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1549]),.i2(intermediate_reg_1[1548]),.o(intermediate_reg_2[774])); 
xor_module xor_module_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1547]),.i2(intermediate_reg_1[1546]),.o(intermediate_reg_2[773])); 
mux_module mux_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1545]),.i2(intermediate_reg_1[1544]),.o(intermediate_reg_2[772]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1543]),.i2(intermediate_reg_1[1542]),.o(intermediate_reg_2[771])); 
mux_module mux_module_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1541]),.i2(intermediate_reg_1[1540]),.o(intermediate_reg_2[770]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1539]),.i2(intermediate_reg_1[1538]),.o(intermediate_reg_2[769]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1537]),.i2(intermediate_reg_1[1536]),.o(intermediate_reg_2[768])); 
mux_module mux_module_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1535]),.i2(intermediate_reg_1[1534]),.o(intermediate_reg_2[767]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1533]),.i2(intermediate_reg_1[1532]),.o(intermediate_reg_2[766]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1531]),.i2(intermediate_reg_1[1530]),.o(intermediate_reg_2[765])); 
xor_module xor_module_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1529]),.i2(intermediate_reg_1[1528]),.o(intermediate_reg_2[764])); 
xor_module xor_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1527]),.i2(intermediate_reg_1[1526]),.o(intermediate_reg_2[763])); 
mux_module mux_module_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1525]),.i2(intermediate_reg_1[1524]),.o(intermediate_reg_2[762]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1523]),.i2(intermediate_reg_1[1522]),.o(intermediate_reg_2[761])); 
mux_module mux_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1521]),.i2(intermediate_reg_1[1520]),.o(intermediate_reg_2[760]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1519]),.i2(intermediate_reg_1[1518]),.o(intermediate_reg_2[759]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1517]),.i2(intermediate_reg_1[1516]),.o(intermediate_reg_2[758]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1515]),.i2(intermediate_reg_1[1514]),.o(intermediate_reg_2[757]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1513]),.i2(intermediate_reg_1[1512]),.o(intermediate_reg_2[756])); 
mux_module mux_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1511]),.i2(intermediate_reg_1[1510]),.o(intermediate_reg_2[755]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1509]),.i2(intermediate_reg_1[1508]),.o(intermediate_reg_2[754])); 
xor_module xor_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1507]),.i2(intermediate_reg_1[1506]),.o(intermediate_reg_2[753])); 
xor_module xor_module_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1505]),.i2(intermediate_reg_1[1504]),.o(intermediate_reg_2[752])); 
xor_module xor_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1503]),.i2(intermediate_reg_1[1502]),.o(intermediate_reg_2[751])); 
xor_module xor_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1501]),.i2(intermediate_reg_1[1500]),.o(intermediate_reg_2[750])); 
xor_module xor_module_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1499]),.i2(intermediate_reg_1[1498]),.o(intermediate_reg_2[749])); 
xor_module xor_module_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1497]),.i2(intermediate_reg_1[1496]),.o(intermediate_reg_2[748])); 
xor_module xor_module_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1495]),.i2(intermediate_reg_1[1494]),.o(intermediate_reg_2[747])); 
xor_module xor_module_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1493]),.i2(intermediate_reg_1[1492]),.o(intermediate_reg_2[746])); 
xor_module xor_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1491]),.i2(intermediate_reg_1[1490]),.o(intermediate_reg_2[745])); 
xor_module xor_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1489]),.i2(intermediate_reg_1[1488]),.o(intermediate_reg_2[744])); 
mux_module mux_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1487]),.i2(intermediate_reg_1[1486]),.o(intermediate_reg_2[743]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1485]),.i2(intermediate_reg_1[1484]),.o(intermediate_reg_2[742]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1483]),.i2(intermediate_reg_1[1482]),.o(intermediate_reg_2[741])); 
xor_module xor_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1481]),.i2(intermediate_reg_1[1480]),.o(intermediate_reg_2[740])); 
mux_module mux_module_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1479]),.i2(intermediate_reg_1[1478]),.o(intermediate_reg_2[739]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1477]),.i2(intermediate_reg_1[1476]),.o(intermediate_reg_2[738]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1475]),.i2(intermediate_reg_1[1474]),.o(intermediate_reg_2[737]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1473]),.i2(intermediate_reg_1[1472]),.o(intermediate_reg_2[736]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1471]),.i2(intermediate_reg_1[1470]),.o(intermediate_reg_2[735])); 
mux_module mux_module_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1469]),.i2(intermediate_reg_1[1468]),.o(intermediate_reg_2[734]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1467]),.i2(intermediate_reg_1[1466]),.o(intermediate_reg_2[733]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1465]),.i2(intermediate_reg_1[1464]),.o(intermediate_reg_2[732])); 
xor_module xor_module_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1463]),.i2(intermediate_reg_1[1462]),.o(intermediate_reg_2[731])); 
mux_module mux_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1461]),.i2(intermediate_reg_1[1460]),.o(intermediate_reg_2[730]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1459]),.i2(intermediate_reg_1[1458]),.o(intermediate_reg_2[729]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1457]),.i2(intermediate_reg_1[1456]),.o(intermediate_reg_2[728])); 
xor_module xor_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1455]),.i2(intermediate_reg_1[1454]),.o(intermediate_reg_2[727])); 
mux_module mux_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1453]),.i2(intermediate_reg_1[1452]),.o(intermediate_reg_2[726]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1451]),.i2(intermediate_reg_1[1450]),.o(intermediate_reg_2[725])); 
xor_module xor_module_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1449]),.i2(intermediate_reg_1[1448]),.o(intermediate_reg_2[724])); 
xor_module xor_module_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1447]),.i2(intermediate_reg_1[1446]),.o(intermediate_reg_2[723])); 
xor_module xor_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1445]),.i2(intermediate_reg_1[1444]),.o(intermediate_reg_2[722])); 
mux_module mux_module_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1443]),.i2(intermediate_reg_1[1442]),.o(intermediate_reg_2[721]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1441]),.i2(intermediate_reg_1[1440]),.o(intermediate_reg_2[720]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1439]),.i2(intermediate_reg_1[1438]),.o(intermediate_reg_2[719])); 
mux_module mux_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1437]),.i2(intermediate_reg_1[1436]),.o(intermediate_reg_2[718]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1435]),.i2(intermediate_reg_1[1434]),.o(intermediate_reg_2[717]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1433]),.i2(intermediate_reg_1[1432]),.o(intermediate_reg_2[716]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1431]),.i2(intermediate_reg_1[1430]),.o(intermediate_reg_2[715])); 
mux_module mux_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1429]),.i2(intermediate_reg_1[1428]),.o(intermediate_reg_2[714]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1427]),.i2(intermediate_reg_1[1426]),.o(intermediate_reg_2[713]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1425]),.i2(intermediate_reg_1[1424]),.o(intermediate_reg_2[712]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1423]),.i2(intermediate_reg_1[1422]),.o(intermediate_reg_2[711]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1421]),.i2(intermediate_reg_1[1420]),.o(intermediate_reg_2[710])); 
mux_module mux_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1419]),.i2(intermediate_reg_1[1418]),.o(intermediate_reg_2[709]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1417]),.i2(intermediate_reg_1[1416]),.o(intermediate_reg_2[708])); 
xor_module xor_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1415]),.i2(intermediate_reg_1[1414]),.o(intermediate_reg_2[707])); 
mux_module mux_module_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1413]),.i2(intermediate_reg_1[1412]),.o(intermediate_reg_2[706]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1411]),.i2(intermediate_reg_1[1410]),.o(intermediate_reg_2[705]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1409]),.i2(intermediate_reg_1[1408]),.o(intermediate_reg_2[704]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1407]),.i2(intermediate_reg_1[1406]),.o(intermediate_reg_2[703]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1405]),.i2(intermediate_reg_1[1404]),.o(intermediate_reg_2[702]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1403]),.i2(intermediate_reg_1[1402]),.o(intermediate_reg_2[701])); 
xor_module xor_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1401]),.i2(intermediate_reg_1[1400]),.o(intermediate_reg_2[700])); 
xor_module xor_module_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1399]),.i2(intermediate_reg_1[1398]),.o(intermediate_reg_2[699])); 
xor_module xor_module_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1397]),.i2(intermediate_reg_1[1396]),.o(intermediate_reg_2[698])); 
mux_module mux_module_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1395]),.i2(intermediate_reg_1[1394]),.o(intermediate_reg_2[697]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1393]),.i2(intermediate_reg_1[1392]),.o(intermediate_reg_2[696])); 
mux_module mux_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1391]),.i2(intermediate_reg_1[1390]),.o(intermediate_reg_2[695]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1389]),.i2(intermediate_reg_1[1388]),.o(intermediate_reg_2[694])); 
mux_module mux_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1387]),.i2(intermediate_reg_1[1386]),.o(intermediate_reg_2[693]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1385]),.i2(intermediate_reg_1[1384]),.o(intermediate_reg_2[692])); 
xor_module xor_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1383]),.i2(intermediate_reg_1[1382]),.o(intermediate_reg_2[691])); 
mux_module mux_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1381]),.i2(intermediate_reg_1[1380]),.o(intermediate_reg_2[690]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1379]),.i2(intermediate_reg_1[1378]),.o(intermediate_reg_2[689])); 
mux_module mux_module_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1377]),.i2(intermediate_reg_1[1376]),.o(intermediate_reg_2[688]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1375]),.i2(intermediate_reg_1[1374]),.o(intermediate_reg_2[687])); 
xor_module xor_module_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1373]),.i2(intermediate_reg_1[1372]),.o(intermediate_reg_2[686])); 
mux_module mux_module_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1371]),.i2(intermediate_reg_1[1370]),.o(intermediate_reg_2[685]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1369]),.i2(intermediate_reg_1[1368]),.o(intermediate_reg_2[684]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1367]),.i2(intermediate_reg_1[1366]),.o(intermediate_reg_2[683])); 
mux_module mux_module_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1365]),.i2(intermediate_reg_1[1364]),.o(intermediate_reg_2[682]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1363]),.i2(intermediate_reg_1[1362]),.o(intermediate_reg_2[681]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1361]),.i2(intermediate_reg_1[1360]),.o(intermediate_reg_2[680]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1359]),.i2(intermediate_reg_1[1358]),.o(intermediate_reg_2[679])); 
mux_module mux_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1357]),.i2(intermediate_reg_1[1356]),.o(intermediate_reg_2[678]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1355]),.i2(intermediate_reg_1[1354]),.o(intermediate_reg_2[677]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1353]),.i2(intermediate_reg_1[1352]),.o(intermediate_reg_2[676])); 
mux_module mux_module_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1351]),.i2(intermediate_reg_1[1350]),.o(intermediate_reg_2[675]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1349]),.i2(intermediate_reg_1[1348]),.o(intermediate_reg_2[674])); 
mux_module mux_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1347]),.i2(intermediate_reg_1[1346]),.o(intermediate_reg_2[673]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1345]),.i2(intermediate_reg_1[1344]),.o(intermediate_reg_2[672]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1343]),.i2(intermediate_reg_1[1342]),.o(intermediate_reg_2[671]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1341]),.i2(intermediate_reg_1[1340]),.o(intermediate_reg_2[670]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1339]),.i2(intermediate_reg_1[1338]),.o(intermediate_reg_2[669])); 
xor_module xor_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1337]),.i2(intermediate_reg_1[1336]),.o(intermediate_reg_2[668])); 
xor_module xor_module_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1335]),.i2(intermediate_reg_1[1334]),.o(intermediate_reg_2[667])); 
mux_module mux_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1333]),.i2(intermediate_reg_1[1332]),.o(intermediate_reg_2[666]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1331]),.i2(intermediate_reg_1[1330]),.o(intermediate_reg_2[665])); 
mux_module mux_module_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1329]),.i2(intermediate_reg_1[1328]),.o(intermediate_reg_2[664]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1327]),.i2(intermediate_reg_1[1326]),.o(intermediate_reg_2[663])); 
mux_module mux_module_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1325]),.i2(intermediate_reg_1[1324]),.o(intermediate_reg_2[662]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1323]),.i2(intermediate_reg_1[1322]),.o(intermediate_reg_2[661]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1321]),.i2(intermediate_reg_1[1320]),.o(intermediate_reg_2[660])); 
mux_module mux_module_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1319]),.i2(intermediate_reg_1[1318]),.o(intermediate_reg_2[659]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1317]),.i2(intermediate_reg_1[1316]),.o(intermediate_reg_2[658]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1315]),.i2(intermediate_reg_1[1314]),.o(intermediate_reg_2[657])); 
xor_module xor_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1313]),.i2(intermediate_reg_1[1312]),.o(intermediate_reg_2[656])); 
mux_module mux_module_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1311]),.i2(intermediate_reg_1[1310]),.o(intermediate_reg_2[655]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1309]),.i2(intermediate_reg_1[1308]),.o(intermediate_reg_2[654]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1307]),.i2(intermediate_reg_1[1306]),.o(intermediate_reg_2[653])); 
mux_module mux_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1305]),.i2(intermediate_reg_1[1304]),.o(intermediate_reg_2[652]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1303]),.i2(intermediate_reg_1[1302]),.o(intermediate_reg_2[651])); 
mux_module mux_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1301]),.i2(intermediate_reg_1[1300]),.o(intermediate_reg_2[650]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1299]),.i2(intermediate_reg_1[1298]),.o(intermediate_reg_2[649])); 
mux_module mux_module_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1297]),.i2(intermediate_reg_1[1296]),.o(intermediate_reg_2[648]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1295]),.i2(intermediate_reg_1[1294]),.o(intermediate_reg_2[647]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1293]),.i2(intermediate_reg_1[1292]),.o(intermediate_reg_2[646]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1291]),.i2(intermediate_reg_1[1290]),.o(intermediate_reg_2[645]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1289]),.i2(intermediate_reg_1[1288]),.o(intermediate_reg_2[644]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1287]),.i2(intermediate_reg_1[1286]),.o(intermediate_reg_2[643]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1285]),.i2(intermediate_reg_1[1284]),.o(intermediate_reg_2[642])); 
xor_module xor_module_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1283]),.i2(intermediate_reg_1[1282]),.o(intermediate_reg_2[641])); 
xor_module xor_module_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1281]),.i2(intermediate_reg_1[1280]),.o(intermediate_reg_2[640])); 
mux_module mux_module_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1279]),.i2(intermediate_reg_1[1278]),.o(intermediate_reg_2[639]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1277]),.i2(intermediate_reg_1[1276]),.o(intermediate_reg_2[638])); 
mux_module mux_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1275]),.i2(intermediate_reg_1[1274]),.o(intermediate_reg_2[637]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1273]),.i2(intermediate_reg_1[1272]),.o(intermediate_reg_2[636]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1271]),.i2(intermediate_reg_1[1270]),.o(intermediate_reg_2[635]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1269]),.i2(intermediate_reg_1[1268]),.o(intermediate_reg_2[634])); 
mux_module mux_module_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1267]),.i2(intermediate_reg_1[1266]),.o(intermediate_reg_2[633]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1265]),.i2(intermediate_reg_1[1264]),.o(intermediate_reg_2[632]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1263]),.i2(intermediate_reg_1[1262]),.o(intermediate_reg_2[631]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1261]),.i2(intermediate_reg_1[1260]),.o(intermediate_reg_2[630])); 
mux_module mux_module_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1259]),.i2(intermediate_reg_1[1258]),.o(intermediate_reg_2[629]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1257]),.i2(intermediate_reg_1[1256]),.o(intermediate_reg_2[628])); 
xor_module xor_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1255]),.i2(intermediate_reg_1[1254]),.o(intermediate_reg_2[627])); 
mux_module mux_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1253]),.i2(intermediate_reg_1[1252]),.o(intermediate_reg_2[626]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1251]),.i2(intermediate_reg_1[1250]),.o(intermediate_reg_2[625])); 
mux_module mux_module_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1249]),.i2(intermediate_reg_1[1248]),.o(intermediate_reg_2[624]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1247]),.i2(intermediate_reg_1[1246]),.o(intermediate_reg_2[623]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1245]),.i2(intermediate_reg_1[1244]),.o(intermediate_reg_2[622]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1243]),.i2(intermediate_reg_1[1242]),.o(intermediate_reg_2[621])); 
mux_module mux_module_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1241]),.i2(intermediate_reg_1[1240]),.o(intermediate_reg_2[620]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1239]),.i2(intermediate_reg_1[1238]),.o(intermediate_reg_2[619]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1237]),.i2(intermediate_reg_1[1236]),.o(intermediate_reg_2[618])); 
xor_module xor_module_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1235]),.i2(intermediate_reg_1[1234]),.o(intermediate_reg_2[617])); 
mux_module mux_module_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1233]),.i2(intermediate_reg_1[1232]),.o(intermediate_reg_2[616]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1231]),.i2(intermediate_reg_1[1230]),.o(intermediate_reg_2[615]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1229]),.i2(intermediate_reg_1[1228]),.o(intermediate_reg_2[614]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1227]),.i2(intermediate_reg_1[1226]),.o(intermediate_reg_2[613]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1225]),.i2(intermediate_reg_1[1224]),.o(intermediate_reg_2[612]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1223]),.i2(intermediate_reg_1[1222]),.o(intermediate_reg_2[611]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1221]),.i2(intermediate_reg_1[1220]),.o(intermediate_reg_2[610])); 
xor_module xor_module_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1219]),.i2(intermediate_reg_1[1218]),.o(intermediate_reg_2[609])); 
xor_module xor_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1217]),.i2(intermediate_reg_1[1216]),.o(intermediate_reg_2[608])); 
mux_module mux_module_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1215]),.i2(intermediate_reg_1[1214]),.o(intermediate_reg_2[607]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1213]),.i2(intermediate_reg_1[1212]),.o(intermediate_reg_2[606]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1211]),.i2(intermediate_reg_1[1210]),.o(intermediate_reg_2[605])); 
mux_module mux_module_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1209]),.i2(intermediate_reg_1[1208]),.o(intermediate_reg_2[604]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1207]),.i2(intermediate_reg_1[1206]),.o(intermediate_reg_2[603]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1205]),.i2(intermediate_reg_1[1204]),.o(intermediate_reg_2[602]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1203]),.i2(intermediate_reg_1[1202]),.o(intermediate_reg_2[601])); 
mux_module mux_module_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1201]),.i2(intermediate_reg_1[1200]),.o(intermediate_reg_2[600]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1199]),.i2(intermediate_reg_1[1198]),.o(intermediate_reg_2[599])); 
mux_module mux_module_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1197]),.i2(intermediate_reg_1[1196]),.o(intermediate_reg_2[598]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1195]),.i2(intermediate_reg_1[1194]),.o(intermediate_reg_2[597])); 
mux_module mux_module_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1193]),.i2(intermediate_reg_1[1192]),.o(intermediate_reg_2[596]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1191]),.i2(intermediate_reg_1[1190]),.o(intermediate_reg_2[595])); 
xor_module xor_module_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1189]),.i2(intermediate_reg_1[1188]),.o(intermediate_reg_2[594])); 
xor_module xor_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1187]),.i2(intermediate_reg_1[1186]),.o(intermediate_reg_2[593])); 
mux_module mux_module_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1185]),.i2(intermediate_reg_1[1184]),.o(intermediate_reg_2[592]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1183]),.i2(intermediate_reg_1[1182]),.o(intermediate_reg_2[591])); 
mux_module mux_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1181]),.i2(intermediate_reg_1[1180]),.o(intermediate_reg_2[590]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1179]),.i2(intermediate_reg_1[1178]),.o(intermediate_reg_2[589])); 
mux_module mux_module_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1177]),.i2(intermediate_reg_1[1176]),.o(intermediate_reg_2[588]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1175]),.i2(intermediate_reg_1[1174]),.o(intermediate_reg_2[587])); 
mux_module mux_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1173]),.i2(intermediate_reg_1[1172]),.o(intermediate_reg_2[586]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1171]),.i2(intermediate_reg_1[1170]),.o(intermediate_reg_2[585])); 
xor_module xor_module_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1169]),.i2(intermediate_reg_1[1168]),.o(intermediate_reg_2[584])); 
mux_module mux_module_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1167]),.i2(intermediate_reg_1[1166]),.o(intermediate_reg_2[583]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1165]),.i2(intermediate_reg_1[1164]),.o(intermediate_reg_2[582]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1163]),.i2(intermediate_reg_1[1162]),.o(intermediate_reg_2[581])); 
mux_module mux_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1161]),.i2(intermediate_reg_1[1160]),.o(intermediate_reg_2[580]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1159]),.i2(intermediate_reg_1[1158]),.o(intermediate_reg_2[579]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1157]),.i2(intermediate_reg_1[1156]),.o(intermediate_reg_2[578]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1155]),.i2(intermediate_reg_1[1154]),.o(intermediate_reg_2[577])); 
xor_module xor_module_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1153]),.i2(intermediate_reg_1[1152]),.o(intermediate_reg_2[576])); 
xor_module xor_module_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1151]),.i2(intermediate_reg_1[1150]),.o(intermediate_reg_2[575])); 
mux_module mux_module_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1149]),.i2(intermediate_reg_1[1148]),.o(intermediate_reg_2[574]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1147]),.i2(intermediate_reg_1[1146]),.o(intermediate_reg_2[573]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1145]),.i2(intermediate_reg_1[1144]),.o(intermediate_reg_2[572])); 
xor_module xor_module_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1143]),.i2(intermediate_reg_1[1142]),.o(intermediate_reg_2[571])); 
xor_module xor_module_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1141]),.i2(intermediate_reg_1[1140]),.o(intermediate_reg_2[570])); 
mux_module mux_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1139]),.i2(intermediate_reg_1[1138]),.o(intermediate_reg_2[569]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1137]),.i2(intermediate_reg_1[1136]),.o(intermediate_reg_2[568])); 
xor_module xor_module_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1135]),.i2(intermediate_reg_1[1134]),.o(intermediate_reg_2[567])); 
xor_module xor_module_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1133]),.i2(intermediate_reg_1[1132]),.o(intermediate_reg_2[566])); 
xor_module xor_module_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1131]),.i2(intermediate_reg_1[1130]),.o(intermediate_reg_2[565])); 
mux_module mux_module_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1129]),.i2(intermediate_reg_1[1128]),.o(intermediate_reg_2[564]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1127]),.i2(intermediate_reg_1[1126]),.o(intermediate_reg_2[563])); 
mux_module mux_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1125]),.i2(intermediate_reg_1[1124]),.o(intermediate_reg_2[562]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1123]),.i2(intermediate_reg_1[1122]),.o(intermediate_reg_2[561])); 
mux_module mux_module_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1121]),.i2(intermediate_reg_1[1120]),.o(intermediate_reg_2[560]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1119]),.i2(intermediate_reg_1[1118]),.o(intermediate_reg_2[559])); 
mux_module mux_module_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1117]),.i2(intermediate_reg_1[1116]),.o(intermediate_reg_2[558]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1115]),.i2(intermediate_reg_1[1114]),.o(intermediate_reg_2[557]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1113]),.i2(intermediate_reg_1[1112]),.o(intermediate_reg_2[556]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1111]),.i2(intermediate_reg_1[1110]),.o(intermediate_reg_2[555]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1109]),.i2(intermediate_reg_1[1108]),.o(intermediate_reg_2[554])); 
mux_module mux_module_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1107]),.i2(intermediate_reg_1[1106]),.o(intermediate_reg_2[553]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1105]),.i2(intermediate_reg_1[1104]),.o(intermediate_reg_2[552]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1103]),.i2(intermediate_reg_1[1102]),.o(intermediate_reg_2[551])); 
xor_module xor_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1101]),.i2(intermediate_reg_1[1100]),.o(intermediate_reg_2[550])); 
xor_module xor_module_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1099]),.i2(intermediate_reg_1[1098]),.o(intermediate_reg_2[549])); 
xor_module xor_module_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1097]),.i2(intermediate_reg_1[1096]),.o(intermediate_reg_2[548])); 
mux_module mux_module_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1095]),.i2(intermediate_reg_1[1094]),.o(intermediate_reg_2[547]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1093]),.i2(intermediate_reg_1[1092]),.o(intermediate_reg_2[546]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1091]),.i2(intermediate_reg_1[1090]),.o(intermediate_reg_2[545]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1089]),.i2(intermediate_reg_1[1088]),.o(intermediate_reg_2[544]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1087]),.i2(intermediate_reg_1[1086]),.o(intermediate_reg_2[543])); 
xor_module xor_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1085]),.i2(intermediate_reg_1[1084]),.o(intermediate_reg_2[542])); 
xor_module xor_module_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1083]),.i2(intermediate_reg_1[1082]),.o(intermediate_reg_2[541])); 
xor_module xor_module_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1081]),.i2(intermediate_reg_1[1080]),.o(intermediate_reg_2[540])); 
xor_module xor_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1079]),.i2(intermediate_reg_1[1078]),.o(intermediate_reg_2[539])); 
mux_module mux_module_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1077]),.i2(intermediate_reg_1[1076]),.o(intermediate_reg_2[538]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1075]),.i2(intermediate_reg_1[1074]),.o(intermediate_reg_2[537]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1073]),.i2(intermediate_reg_1[1072]),.o(intermediate_reg_2[536])); 
mux_module mux_module_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1071]),.i2(intermediate_reg_1[1070]),.o(intermediate_reg_2[535]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1069]),.i2(intermediate_reg_1[1068]),.o(intermediate_reg_2[534]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1067]),.i2(intermediate_reg_1[1066]),.o(intermediate_reg_2[533]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1065]),.i2(intermediate_reg_1[1064]),.o(intermediate_reg_2[532])); 
mux_module mux_module_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1063]),.i2(intermediate_reg_1[1062]),.o(intermediate_reg_2[531]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1061]),.i2(intermediate_reg_1[1060]),.o(intermediate_reg_2[530])); 
xor_module xor_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1059]),.i2(intermediate_reg_1[1058]),.o(intermediate_reg_2[529])); 
mux_module mux_module_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1057]),.i2(intermediate_reg_1[1056]),.o(intermediate_reg_2[528]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1055]),.i2(intermediate_reg_1[1054]),.o(intermediate_reg_2[527]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1053]),.i2(intermediate_reg_1[1052]),.o(intermediate_reg_2[526]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1051]),.i2(intermediate_reg_1[1050]),.o(intermediate_reg_2[525])); 
xor_module xor_module_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1049]),.i2(intermediate_reg_1[1048]),.o(intermediate_reg_2[524])); 
mux_module mux_module_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1047]),.i2(intermediate_reg_1[1046]),.o(intermediate_reg_2[523]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1045]),.i2(intermediate_reg_1[1044]),.o(intermediate_reg_2[522])); 
mux_module mux_module_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1043]),.i2(intermediate_reg_1[1042]),.o(intermediate_reg_2[521]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1041]),.i2(intermediate_reg_1[1040]),.o(intermediate_reg_2[520])); 
xor_module xor_module_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1039]),.i2(intermediate_reg_1[1038]),.o(intermediate_reg_2[519])); 
xor_module xor_module_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1037]),.i2(intermediate_reg_1[1036]),.o(intermediate_reg_2[518])); 
mux_module mux_module_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1035]),.i2(intermediate_reg_1[1034]),.o(intermediate_reg_2[517]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1033]),.i2(intermediate_reg_1[1032]),.o(intermediate_reg_2[516]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1031]),.i2(intermediate_reg_1[1030]),.o(intermediate_reg_2[515]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1029]),.i2(intermediate_reg_1[1028]),.o(intermediate_reg_2[514])); 
xor_module xor_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513])); 
mux_module mux_module_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509])); 
mux_module mux_module_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507])); 
xor_module xor_module_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506])); 
xor_module xor_module_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505])); 
mux_module mux_module_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503])); 
mux_module mux_module_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498])); 
mux_module mux_module_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494])); 
mux_module mux_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492])); 
mux_module mux_module_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488])); 
xor_module xor_module_inst_2_516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487])); 
xor_module xor_module_inst_2_517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486])); 
xor_module xor_module_inst_2_518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485])); 
xor_module xor_module_inst_2_519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484])); 
mux_module mux_module_inst_2_520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482])); 
xor_module xor_module_inst_2_522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481])); 
mux_module mux_module_inst_2_523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
xor_module xor_module_inst_2_525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478])); 
mux_module mux_module_inst_2_526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476])); 
mux_module mux_module_inst_2_528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474])); 
xor_module xor_module_inst_2_530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473])); 
mux_module mux_module_inst_2_531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470])); 
mux_module mux_module_inst_2_534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466])); 
xor_module xor_module_inst_2_538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465])); 
mux_module mux_module_inst_2_539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458])); 
xor_module xor_module_inst_2_546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457])); 
xor_module xor_module_inst_2_547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456])); 
xor_module xor_module_inst_2_548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455])); 
xor_module xor_module_inst_2_549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454])); 
xor_module xor_module_inst_2_550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453])); 
mux_module mux_module_inst_2_551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450])); 
mux_module mux_module_inst_2_554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448])); 
xor_module xor_module_inst_2_556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447])); 
mux_module mux_module_inst_2_557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445])); 
mux_module mux_module_inst_2_559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_560(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443])); 
xor_module xor_module_inst_2_561(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442])); 
xor_module xor_module_inst_2_562(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441])); 
xor_module xor_module_inst_2_563(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440])); 
mux_module mux_module_inst_2_564(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_565(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438])); 
mux_module mux_module_inst_2_566(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_567(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436])); 
xor_module xor_module_inst_2_568(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435])); 
mux_module mux_module_inst_2_569(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_570(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_571(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432])); 
mux_module mux_module_inst_2_572(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_573(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430])); 
xor_module xor_module_inst_2_574(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429])); 
xor_module xor_module_inst_2_575(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428])); 
xor_module xor_module_inst_2_576(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427])); 
mux_module mux_module_inst_2_577(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_578(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425])); 
mux_module mux_module_inst_2_579(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_580(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_581(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_582(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_583(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420])); 
mux_module mux_module_inst_2_584(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_585(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418])); 
mux_module mux_module_inst_2_586(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_587(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416])); 
mux_module mux_module_inst_2_588(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_589(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_590(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413])); 
mux_module mux_module_inst_2_591(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_592(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411])); 
xor_module xor_module_inst_2_593(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410])); 
mux_module mux_module_inst_2_594(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_595(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_596(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407])); 
xor_module xor_module_inst_2_597(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406])); 
mux_module mux_module_inst_2_598(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_599(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404])); 
xor_module xor_module_inst_2_600(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403])); 
mux_module mux_module_inst_2_601(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_602(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401])); 
xor_module xor_module_inst_2_603(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400])); 
xor_module xor_module_inst_2_604(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399])); 
mux_module mux_module_inst_2_605(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_606(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_607(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396])); 
xor_module xor_module_inst_2_608(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395])); 
xor_module xor_module_inst_2_609(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394])); 
xor_module xor_module_inst_2_610(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393])); 
xor_module xor_module_inst_2_611(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392])); 
xor_module xor_module_inst_2_612(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391])); 
xor_module xor_module_inst_2_613(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390])); 
mux_module mux_module_inst_2_614(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_615(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_616(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_617(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_618(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_619(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_620(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383])); 
xor_module xor_module_inst_2_621(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382])); 
xor_module xor_module_inst_2_622(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
xor_module xor_module_inst_2_623(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
mux_module mux_module_inst_2_624(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_625(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378])); 
xor_module xor_module_inst_2_626(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377])); 
mux_module mux_module_inst_2_627(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_628(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_629(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_630(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373])); 
xor_module xor_module_inst_2_631(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372])); 
xor_module xor_module_inst_2_632(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371])); 
xor_module xor_module_inst_2_633(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
mux_module mux_module_inst_2_634(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_635(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368])); 
xor_module xor_module_inst_2_636(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367])); 
xor_module xor_module_inst_2_637(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366])); 
xor_module xor_module_inst_2_638(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365])); 
xor_module xor_module_inst_2_639(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
xor_module xor_module_inst_2_640(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363])); 
xor_module xor_module_inst_2_641(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362])); 
mux_module mux_module_inst_2_642(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_643(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_644(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_645(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
mux_module mux_module_inst_2_646(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_647(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356])); 
mux_module mux_module_inst_2_648(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_649(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354])); 
xor_module xor_module_inst_2_650(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353])); 
mux_module mux_module_inst_2_651(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_652(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351])); 
xor_module xor_module_inst_2_653(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350])); 
mux_module mux_module_inst_2_654(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_655(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_656(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
mux_module mux_module_inst_2_657(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_658(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_659(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_660(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_661(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342])); 
xor_module xor_module_inst_2_662(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341])); 
xor_module xor_module_inst_2_663(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340])); 
mux_module mux_module_inst_2_664(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_665(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_666(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_667(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_668(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_669(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334])); 
xor_module xor_module_inst_2_670(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333])); 
xor_module xor_module_inst_2_671(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332])); 
xor_module xor_module_inst_2_672(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331])); 
xor_module xor_module_inst_2_673(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
mux_module mux_module_inst_2_674(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_675(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_676(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
xor_module xor_module_inst_2_677(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326])); 
mux_module mux_module_inst_2_678(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_679(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_680(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323])); 
mux_module mux_module_inst_2_681(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_682(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_683(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
mux_module mux_module_inst_2_684(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_685(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318])); 
mux_module mux_module_inst_2_686(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_687(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316])); 
mux_module mux_module_inst_2_688(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_689(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314])); 
mux_module mux_module_inst_2_690(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_691(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312])); 
mux_module mux_module_inst_2_692(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_693(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_694(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309])); 
xor_module xor_module_inst_2_695(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308])); 
xor_module xor_module_inst_2_696(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307])); 
xor_module xor_module_inst_2_697(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306])); 
xor_module xor_module_inst_2_698(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305])); 
mux_module mux_module_inst_2_699(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_700(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
mux_module mux_module_inst_2_701(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_702(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_703(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300])); 
mux_module mux_module_inst_2_704(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_705(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298])); 
mux_module mux_module_inst_2_706(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_707(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
mux_module mux_module_inst_2_708(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_709(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294])); 
mux_module mux_module_inst_2_710(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_711(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292])); 
mux_module mux_module_inst_2_712(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_713(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_714(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_715(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288])); 
mux_module mux_module_inst_2_716(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_717(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_718(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
xor_module xor_module_inst_2_719(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284])); 
xor_module xor_module_inst_2_720(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
xor_module xor_module_inst_2_721(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282])); 
mux_module mux_module_inst_2_722(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_723(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_724(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279])); 
xor_module xor_module_inst_2_725(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278])); 
mux_module mux_module_inst_2_726(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_727(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_728(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_729(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
mux_module mux_module_inst_2_730(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_731(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
xor_module xor_module_inst_2_732(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
mux_module mux_module_inst_2_733(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_734(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_735(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_736(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_737(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_738(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_739(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_740(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_741(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_742(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_743(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
xor_module xor_module_inst_2_744(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259])); 
mux_module mux_module_inst_2_745(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_746(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_747(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
xor_module xor_module_inst_2_748(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255])); 
mux_module mux_module_inst_2_749(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_750(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_751(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_752(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_753(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_754(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_755(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248])); 
xor_module xor_module_inst_2_756(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247])); 
mux_module mux_module_inst_2_757(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_758(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
xor_module xor_module_inst_2_759(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244])); 
mux_module mux_module_inst_2_760(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_761(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242])); 
xor_module xor_module_inst_2_762(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
mux_module mux_module_inst_2_763(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_764(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239])); 
mux_module mux_module_inst_2_765(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_766(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
mux_module mux_module_inst_2_767(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_768(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235])); 
xor_module xor_module_inst_2_769(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
mux_module mux_module_inst_2_770(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_771(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_772(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_773(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_774(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229])); 
xor_module xor_module_inst_2_775(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
xor_module xor_module_inst_2_776(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227])); 
xor_module xor_module_inst_2_777(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
xor_module xor_module_inst_2_778(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
xor_module xor_module_inst_2_779(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224])); 
mux_module mux_module_inst_2_780(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_781(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
mux_module mux_module_inst_2_782(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_783(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_784(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_785(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
mux_module mux_module_inst_2_786(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_787(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216])); 
mux_module mux_module_inst_2_788(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_789(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_790(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
xor_module xor_module_inst_2_791(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
xor_module xor_module_inst_2_792(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
xor_module xor_module_inst_2_793(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
mux_module mux_module_inst_2_794(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_795(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208])); 
mux_module mux_module_inst_2_796(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_797(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
xor_module xor_module_inst_2_798(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
mux_module mux_module_inst_2_799(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_800(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203])); 
xor_module xor_module_inst_2_801(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202])); 
mux_module mux_module_inst_2_802(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_803(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200])); 
xor_module xor_module_inst_2_804(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
mux_module mux_module_inst_2_805(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_806(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_807(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
xor_module xor_module_inst_2_808(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195])); 
xor_module xor_module_inst_2_809(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194])); 
mux_module mux_module_inst_2_810(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_811(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
xor_module xor_module_inst_2_812(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
mux_module mux_module_inst_2_813(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_814(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_815(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
xor_module xor_module_inst_2_816(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
xor_module xor_module_inst_2_817(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186])); 
xor_module xor_module_inst_2_818(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185])); 
xor_module xor_module_inst_2_819(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
mux_module mux_module_inst_2_820(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_821(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_822(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_823(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_824(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_825(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_826(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_827(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_828(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_829(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174])); 
xor_module xor_module_inst_2_830(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
mux_module mux_module_inst_2_831(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_832(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
xor_module xor_module_inst_2_833(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
xor_module xor_module_inst_2_834(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169])); 
mux_module mux_module_inst_2_835(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_836(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_837(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_838(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
mux_module mux_module_inst_2_839(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_840(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_841(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_842(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_843(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_844(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_845(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_846(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_847(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_848(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_849(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_850(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153])); 
mux_module mux_module_inst_2_851(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_852(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151])); 
mux_module mux_module_inst_2_853(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_854(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
xor_module xor_module_inst_2_855(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148])); 
mux_module mux_module_inst_2_856(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_857(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_858(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_859(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_860(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_861(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142])); 
mux_module mux_module_inst_2_862(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_863(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140])); 
xor_module xor_module_inst_2_864(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139])); 
xor_module xor_module_inst_2_865(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138])); 
mux_module mux_module_inst_2_866(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_867(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136])); 
mux_module mux_module_inst_2_868(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_869(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_870(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_871(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_872(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131])); 
mux_module mux_module_inst_2_873(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_874(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129])); 
xor_module xor_module_inst_2_875(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
mux_module mux_module_inst_2_876(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_877(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126])); 
mux_module mux_module_inst_2_878(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_879(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_880(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123])); 
mux_module mux_module_inst_2_881(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_882(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_883(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_884(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119])); 
mux_module mux_module_inst_2_885(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_886(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_887(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116])); 
mux_module mux_module_inst_2_888(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_889(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_890(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_891(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_892(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111])); 
xor_module xor_module_inst_2_893(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
xor_module xor_module_inst_2_894(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
mux_module mux_module_inst_2_895(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_896(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107])); 
xor_module xor_module_inst_2_897(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
mux_module mux_module_inst_2_898(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_899(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_900(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
mux_module mux_module_inst_2_901(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_902(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_903(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_904(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99])); 
mux_module mux_module_inst_2_905(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_906(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_907(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_908(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_909(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94])); 
mux_module mux_module_inst_2_910(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_911(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92])); 
xor_module xor_module_inst_2_912(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91])); 
mux_module mux_module_inst_2_913(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_914(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89])); 
mux_module mux_module_inst_2_915(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_916(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
mux_module mux_module_inst_2_917(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_918(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_919(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
xor_module xor_module_inst_2_920(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
mux_module mux_module_inst_2_921(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_922(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
mux_module mux_module_inst_2_923(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_924(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79])); 
mux_module mux_module_inst_2_925(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_926(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_927(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76])); 
xor_module xor_module_inst_2_928(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
xor_module xor_module_inst_2_929(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74])); 
mux_module mux_module_inst_2_930(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_931(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_932(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71])); 
xor_module xor_module_inst_2_933(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
xor_module xor_module_inst_2_934(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69])); 
xor_module xor_module_inst_2_935(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68])); 
mux_module mux_module_inst_2_936(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_937(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66])); 
xor_module xor_module_inst_2_938(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65])); 
mux_module mux_module_inst_2_939(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_940(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
xor_module xor_module_inst_2_941(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
mux_module mux_module_inst_2_942(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_943(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_944(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_945(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
xor_module xor_module_inst_2_946(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57])); 
mux_module mux_module_inst_2_947(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_948(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55])); 
xor_module xor_module_inst_2_949(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54])); 
xor_module xor_module_inst_2_950(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
xor_module xor_module_inst_2_951(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
xor_module xor_module_inst_2_952(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51])); 
xor_module xor_module_inst_2_953(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
xor_module xor_module_inst_2_954(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
xor_module xor_module_inst_2_955(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48])); 
mux_module mux_module_inst_2_956(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_957(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_958(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45])); 
mux_module mux_module_inst_2_959(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_960(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_961(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_962(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_963(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_964(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39])); 
mux_module mux_module_inst_2_965(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_966(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
mux_module mux_module_inst_2_967(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_968(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35])); 
mux_module mux_module_inst_2_969(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_970(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_971(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_972(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
xor_module xor_module_inst_2_973(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
mux_module mux_module_inst_2_974(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_975(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
xor_module xor_module_inst_2_976(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27])); 
xor_module xor_module_inst_2_977(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26])); 
xor_module xor_module_inst_2_978(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25])); 
mux_module mux_module_inst_2_979(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_980(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23])); 
mux_module mux_module_inst_2_981(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_982(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21])); 
xor_module xor_module_inst_2_983(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20])); 
xor_module xor_module_inst_2_984(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
xor_module xor_module_inst_2_985(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18])); 
xor_module xor_module_inst_2_986(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17])); 
xor_module xor_module_inst_2_987(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
mux_module mux_module_inst_2_988(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_989(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_990(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13])); 
mux_module mux_module_inst_2_991(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_992(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11])); 
mux_module mux_module_inst_2_993(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_994(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
mux_module mux_module_inst_2_995(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_996(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
mux_module mux_module_inst_2_997(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_998(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5])); 
xor_module xor_module_inst_2_999(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
xor_module xor_module_inst_2_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
mux_module mux_module_inst_2_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0]),.sel(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [1003:0] <= intermediate_reg_2; 
outp[1535:1004] <= intermediate_reg_2[531:0] ; 
end 
endmodule 
 

module interface_7(input [1663:0] inp, output reg [3179:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[1663:0] <= inp ; 
outp[3179:1664] <= inp[1515:0] ; 
end 
endmodule 

module interface_8(input [191:0] inp, output reg [529:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[191:0] <= inp ; 
outp[383:192] <= inp ; 
outp[529:384] <= inp[145:0] ; 
end 
endmodule 

module interface_10(input [2623:0] inp, output reg [1055:0] outp, input clk, input reset);
reg [2623:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1311:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308])); 
xor_module xor_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304])); 
xor_module xor_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276])); 
xor_module xor_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271])); 
xor_module xor_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267])); 
xor_module xor_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263])); 
xor_module xor_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255])); 
xor_module xor_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246])); 
xor_module xor_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235])); 
xor_module xor_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234])); 
xor_module xor_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233])); 
xor_module xor_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231])); 
mux_module mux_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
mux_module mux_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209])); 
xor_module xor_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195])); 
mux_module mux_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193])); 
xor_module xor_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190])); 
xor_module xor_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180])); 
xor_module xor_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179])); 
mux_module mux_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169])); 
mux_module mux_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161])); 
mux_module mux_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159])); 
xor_module xor_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154])); 
mux_module mux_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
mux_module mux_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146])); 
xor_module xor_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133])); 
mux_module mux_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
mux_module mux_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122])); 
xor_module xor_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109])); 
mux_module mux_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
xor_module xor_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
xor_module xor_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102])); 
xor_module xor_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
mux_module mux_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095])); 
mux_module mux_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072])); 
mux_module mux_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068])); 
xor_module xor_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
xor_module xor_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059])); 
xor_module xor_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048])); 
xor_module xor_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
xor_module xor_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
xor_module xor_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033])); 
xor_module xor_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
xor_module xor_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
xor_module xor_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022])); 
mux_module mux_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
mux_module mux_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013])); 
mux_module mux_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009])); 
xor_module xor_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
xor_module xor_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
mux_module mux_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001])); 
xor_module xor_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
mux_module mux_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
xor_module xor_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
mux_module mux_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
mux_module mux_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
xor_module xor_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
mux_module mux_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
mux_module mux_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
xor_module xor_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
mux_module mux_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
mux_module mux_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950])); 
mux_module mux_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
xor_module xor_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
xor_module xor_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
xor_module xor_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
xor_module xor_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
mux_module mux_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
mux_module mux_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
xor_module xor_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
mux_module mux_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
xor_module xor_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
xor_module xor_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
xor_module xor_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
xor_module xor_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
xor_module xor_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
xor_module xor_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
xor_module xor_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
mux_module mux_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
mux_module mux_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
mux_module mux_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
mux_module mux_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
mux_module mux_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
xor_module xor_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
xor_module xor_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
xor_module xor_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
xor_module xor_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
mux_module mux_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
xor_module xor_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
xor_module xor_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
xor_module xor_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
mux_module mux_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
mux_module mux_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
mux_module mux_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
mux_module mux_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
mux_module mux_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
xor_module xor_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
xor_module xor_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
xor_module xor_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
mux_module mux_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
mux_module mux_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
xor_module xor_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
xor_module xor_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
mux_module mux_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
xor_module xor_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
xor_module xor_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
xor_module xor_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
xor_module xor_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
xor_module xor_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
xor_module xor_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
xor_module xor_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
xor_module xor_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
mux_module mux_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
xor_module xor_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
xor_module xor_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
mux_module mux_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
xor_module xor_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
xor_module xor_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
xor_module xor_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
xor_module xor_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
xor_module xor_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
mux_module mux_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
xor_module xor_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
mux_module mux_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
xor_module xor_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
mux_module mux_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
mux_module mux_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
xor_module xor_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
mux_module mux_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
mux_module mux_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
xor_module xor_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
xor_module xor_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
xor_module xor_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
xor_module xor_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
mux_module mux_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
mux_module mux_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
xor_module xor_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
xor_module xor_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
xor_module xor_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
xor_module xor_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
xor_module xor_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
mux_module mux_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
mux_module mux_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
xor_module xor_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
xor_module xor_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
xor_module xor_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
xor_module xor_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
mux_module mux_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
xor_module xor_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
xor_module xor_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
xor_module xor_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
xor_module xor_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
mux_module mux_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
xor_module xor_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
mux_module mux_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
xor_module xor_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
mux_module mux_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
mux_module mux_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
mux_module mux_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
mux_module mux_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
mux_module mux_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
xor_module xor_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
xor_module xor_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
xor_module xor_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
xor_module xor_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
mux_module mux_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
xor_module xor_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
mux_module mux_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
xor_module xor_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
xor_module xor_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
mux_module mux_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
xor_module xor_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
mux_module mux_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
mux_module mux_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
xor_module xor_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
mux_module mux_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
xor_module xor_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
xor_module xor_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
mux_module mux_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
xor_module xor_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
xor_module xor_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
xor_module xor_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
mux_module mux_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
xor_module xor_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
mux_module mux_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
mux_module mux_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
mux_module mux_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
mux_module mux_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
xor_module xor_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
xor_module xor_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
mux_module mux_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
mux_module mux_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
mux_module mux_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
xor_module xor_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
xor_module xor_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
xor_module xor_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
xor_module xor_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
xor_module xor_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
xor_module xor_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
mux_module mux_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
xor_module xor_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
mux_module mux_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
xor_module xor_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
mux_module mux_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
mux_module mux_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
mux_module mux_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
mux_module mux_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
mux_module mux_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
mux_module mux_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
mux_module mux_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
xor_module xor_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
mux_module mux_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
xor_module xor_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
xor_module xor_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
mux_module mux_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
xor_module xor_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
xor_module xor_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
xor_module xor_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
xor_module xor_module_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
xor_module xor_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
mux_module mux_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
mux_module mux_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
mux_module mux_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
mux_module mux_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
mux_module mux_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
mux_module mux_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
mux_module mux_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
xor_module xor_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
xor_module xor_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
xor_module xor_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
xor_module xor_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
xor_module xor_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
mux_module mux_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
xor_module xor_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
xor_module xor_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
mux_module mux_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
mux_module mux_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
xor_module xor_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
xor_module xor_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
xor_module xor_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
mux_module mux_module_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
xor_module xor_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
xor_module xor_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
mux_module mux_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
mux_module mux_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
xor_module xor_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
xor_module xor_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
mux_module mux_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
mux_module mux_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
xor_module xor_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
xor_module xor_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
mux_module mux_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
xor_module xor_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
mux_module mux_module_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
mux_module mux_module_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
xor_module xor_module_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
xor_module xor_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
xor_module xor_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
xor_module xor_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
xor_module xor_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
xor_module xor_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
xor_module xor_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
mux_module mux_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
xor_module xor_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
mux_module mux_module_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
mux_module mux_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
mux_module mux_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
mux_module mux_module_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
mux_module mux_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
xor_module xor_module_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
xor_module xor_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
mux_module mux_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
xor_module xor_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
xor_module xor_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
mux_module mux_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
mux_module mux_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
mux_module mux_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
xor_module xor_module_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
xor_module xor_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
xor_module xor_module_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
xor_module xor_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
xor_module xor_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
xor_module xor_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
mux_module mux_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
mux_module mux_module_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
mux_module mux_module_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
mux_module mux_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
xor_module xor_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
xor_module xor_module_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
mux_module mux_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
mux_module mux_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
xor_module xor_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
xor_module xor_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
mux_module mux_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
mux_module mux_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
mux_module mux_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
mux_module mux_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
xor_module xor_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
xor_module xor_module_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
mux_module mux_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
mux_module mux_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
xor_module xor_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
xor_module xor_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
mux_module mux_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
mux_module mux_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
xor_module xor_module_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
xor_module xor_module_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
xor_module xor_module_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
xor_module xor_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
mux_module mux_module_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
mux_module mux_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
mux_module mux_module_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
mux_module mux_module_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
xor_module xor_module_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
xor_module xor_module_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
mux_module mux_module_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
xor_module xor_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
xor_module xor_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
mux_module mux_module_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
mux_module mux_module_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
xor_module xor_module_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
xor_module xor_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
xor_module xor_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
mux_module mux_module_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
mux_module mux_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
mux_module mux_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
mux_module mux_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
mux_module mux_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
mux_module mux_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
mux_module mux_module_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
xor_module xor_module_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
mux_module mux_module_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
mux_module mux_module_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
xor_module xor_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
mux_module mux_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
mux_module mux_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
xor_module xor_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
mux_module mux_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
xor_module xor_module_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
xor_module xor_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
xor_module xor_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
mux_module mux_module_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
xor_module xor_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
mux_module mux_module_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
xor_module xor_module_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
xor_module xor_module_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
xor_module xor_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
mux_module mux_module_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
mux_module mux_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
xor_module xor_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
xor_module xor_module_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
xor_module xor_module_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
mux_module mux_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
xor_module xor_module_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
mux_module mux_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
mux_module mux_module_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
mux_module mux_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
mux_module mux_module_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
xor_module xor_module_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
xor_module xor_module_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
mux_module mux_module_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
xor_module xor_module_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
mux_module mux_module_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
mux_module mux_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
xor_module xor_module_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
mux_module mux_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
mux_module mux_module_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
xor_module xor_module_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
mux_module mux_module_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
mux_module mux_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
mux_module mux_module_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
xor_module xor_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
mux_module mux_module_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
xor_module xor_module_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
mux_module mux_module_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
reg [655:0]intermediate_reg_2; 
 
xor_module xor_module_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1311]),.i2(intermediate_reg_1[1310]),.o(intermediate_reg_2[655])); 
mux_module mux_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1309]),.i2(intermediate_reg_1[1308]),.o(intermediate_reg_2[654]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1307]),.i2(intermediate_reg_1[1306]),.o(intermediate_reg_2[653])); 
xor_module xor_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1305]),.i2(intermediate_reg_1[1304]),.o(intermediate_reg_2[652])); 
mux_module mux_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1303]),.i2(intermediate_reg_1[1302]),.o(intermediate_reg_2[651]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1301]),.i2(intermediate_reg_1[1300]),.o(intermediate_reg_2[650]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1299]),.i2(intermediate_reg_1[1298]),.o(intermediate_reg_2[649]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1297]),.i2(intermediate_reg_1[1296]),.o(intermediate_reg_2[648])); 
xor_module xor_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1295]),.i2(intermediate_reg_1[1294]),.o(intermediate_reg_2[647])); 
mux_module mux_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1293]),.i2(intermediate_reg_1[1292]),.o(intermediate_reg_2[646]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1291]),.i2(intermediate_reg_1[1290]),.o(intermediate_reg_2[645])); 
xor_module xor_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1289]),.i2(intermediate_reg_1[1288]),.o(intermediate_reg_2[644])); 
mux_module mux_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1287]),.i2(intermediate_reg_1[1286]),.o(intermediate_reg_2[643]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1285]),.i2(intermediate_reg_1[1284]),.o(intermediate_reg_2[642])); 
xor_module xor_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1283]),.i2(intermediate_reg_1[1282]),.o(intermediate_reg_2[641])); 
xor_module xor_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1281]),.i2(intermediate_reg_1[1280]),.o(intermediate_reg_2[640])); 
xor_module xor_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1279]),.i2(intermediate_reg_1[1278]),.o(intermediate_reg_2[639])); 
xor_module xor_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1277]),.i2(intermediate_reg_1[1276]),.o(intermediate_reg_2[638])); 
xor_module xor_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1275]),.i2(intermediate_reg_1[1274]),.o(intermediate_reg_2[637])); 
mux_module mux_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1273]),.i2(intermediate_reg_1[1272]),.o(intermediate_reg_2[636]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1271]),.i2(intermediate_reg_1[1270]),.o(intermediate_reg_2[635])); 
mux_module mux_module_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1269]),.i2(intermediate_reg_1[1268]),.o(intermediate_reg_2[634]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1267]),.i2(intermediate_reg_1[1266]),.o(intermediate_reg_2[633]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1265]),.i2(intermediate_reg_1[1264]),.o(intermediate_reg_2[632])); 
xor_module xor_module_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1263]),.i2(intermediate_reg_1[1262]),.o(intermediate_reg_2[631])); 
mux_module mux_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1261]),.i2(intermediate_reg_1[1260]),.o(intermediate_reg_2[630]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1259]),.i2(intermediate_reg_1[1258]),.o(intermediate_reg_2[629])); 
xor_module xor_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1257]),.i2(intermediate_reg_1[1256]),.o(intermediate_reg_2[628])); 
xor_module xor_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1255]),.i2(intermediate_reg_1[1254]),.o(intermediate_reg_2[627])); 
mux_module mux_module_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1253]),.i2(intermediate_reg_1[1252]),.o(intermediate_reg_2[626]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1251]),.i2(intermediate_reg_1[1250]),.o(intermediate_reg_2[625])); 
mux_module mux_module_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1249]),.i2(intermediate_reg_1[1248]),.o(intermediate_reg_2[624]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1247]),.i2(intermediate_reg_1[1246]),.o(intermediate_reg_2[623])); 
mux_module mux_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1245]),.i2(intermediate_reg_1[1244]),.o(intermediate_reg_2[622]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1243]),.i2(intermediate_reg_1[1242]),.o(intermediate_reg_2[621])); 
xor_module xor_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1241]),.i2(intermediate_reg_1[1240]),.o(intermediate_reg_2[620])); 
xor_module xor_module_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1239]),.i2(intermediate_reg_1[1238]),.o(intermediate_reg_2[619])); 
xor_module xor_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1237]),.i2(intermediate_reg_1[1236]),.o(intermediate_reg_2[618])); 
xor_module xor_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1235]),.i2(intermediate_reg_1[1234]),.o(intermediate_reg_2[617])); 
mux_module mux_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1233]),.i2(intermediate_reg_1[1232]),.o(intermediate_reg_2[616]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1231]),.i2(intermediate_reg_1[1230]),.o(intermediate_reg_2[615])); 
mux_module mux_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1229]),.i2(intermediate_reg_1[1228]),.o(intermediate_reg_2[614]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1227]),.i2(intermediate_reg_1[1226]),.o(intermediate_reg_2[613])); 
mux_module mux_module_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1225]),.i2(intermediate_reg_1[1224]),.o(intermediate_reg_2[612]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1223]),.i2(intermediate_reg_1[1222]),.o(intermediate_reg_2[611])); 
xor_module xor_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1221]),.i2(intermediate_reg_1[1220]),.o(intermediate_reg_2[610])); 
mux_module mux_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1219]),.i2(intermediate_reg_1[1218]),.o(intermediate_reg_2[609]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1217]),.i2(intermediate_reg_1[1216]),.o(intermediate_reg_2[608])); 
xor_module xor_module_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1215]),.i2(intermediate_reg_1[1214]),.o(intermediate_reg_2[607])); 
xor_module xor_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1213]),.i2(intermediate_reg_1[1212]),.o(intermediate_reg_2[606])); 
mux_module mux_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1211]),.i2(intermediate_reg_1[1210]),.o(intermediate_reg_2[605]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1209]),.i2(intermediate_reg_1[1208]),.o(intermediate_reg_2[604]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1207]),.i2(intermediate_reg_1[1206]),.o(intermediate_reg_2[603]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1205]),.i2(intermediate_reg_1[1204]),.o(intermediate_reg_2[602])); 
xor_module xor_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1203]),.i2(intermediate_reg_1[1202]),.o(intermediate_reg_2[601])); 
xor_module xor_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1201]),.i2(intermediate_reg_1[1200]),.o(intermediate_reg_2[600])); 
xor_module xor_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1199]),.i2(intermediate_reg_1[1198]),.o(intermediate_reg_2[599])); 
mux_module mux_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1197]),.i2(intermediate_reg_1[1196]),.o(intermediate_reg_2[598]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1195]),.i2(intermediate_reg_1[1194]),.o(intermediate_reg_2[597]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1193]),.i2(intermediate_reg_1[1192]),.o(intermediate_reg_2[596])); 
xor_module xor_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1191]),.i2(intermediate_reg_1[1190]),.o(intermediate_reg_2[595])); 
mux_module mux_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1189]),.i2(intermediate_reg_1[1188]),.o(intermediate_reg_2[594]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1187]),.i2(intermediate_reg_1[1186]),.o(intermediate_reg_2[593]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1185]),.i2(intermediate_reg_1[1184]),.o(intermediate_reg_2[592])); 
xor_module xor_module_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1183]),.i2(intermediate_reg_1[1182]),.o(intermediate_reg_2[591])); 
xor_module xor_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1181]),.i2(intermediate_reg_1[1180]),.o(intermediate_reg_2[590])); 
xor_module xor_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1179]),.i2(intermediate_reg_1[1178]),.o(intermediate_reg_2[589])); 
mux_module mux_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1177]),.i2(intermediate_reg_1[1176]),.o(intermediate_reg_2[588]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1175]),.i2(intermediate_reg_1[1174]),.o(intermediate_reg_2[587])); 
xor_module xor_module_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1173]),.i2(intermediate_reg_1[1172]),.o(intermediate_reg_2[586])); 
mux_module mux_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1171]),.i2(intermediate_reg_1[1170]),.o(intermediate_reg_2[585]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1169]),.i2(intermediate_reg_1[1168]),.o(intermediate_reg_2[584]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1167]),.i2(intermediate_reg_1[1166]),.o(intermediate_reg_2[583]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1165]),.i2(intermediate_reg_1[1164]),.o(intermediate_reg_2[582])); 
xor_module xor_module_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1163]),.i2(intermediate_reg_1[1162]),.o(intermediate_reg_2[581])); 
mux_module mux_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1161]),.i2(intermediate_reg_1[1160]),.o(intermediate_reg_2[580]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1159]),.i2(intermediate_reg_1[1158]),.o(intermediate_reg_2[579])); 
xor_module xor_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1157]),.i2(intermediate_reg_1[1156]),.o(intermediate_reg_2[578])); 
xor_module xor_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1155]),.i2(intermediate_reg_1[1154]),.o(intermediate_reg_2[577])); 
mux_module mux_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1153]),.i2(intermediate_reg_1[1152]),.o(intermediate_reg_2[576]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1151]),.i2(intermediate_reg_1[1150]),.o(intermediate_reg_2[575]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1149]),.i2(intermediate_reg_1[1148]),.o(intermediate_reg_2[574]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1147]),.i2(intermediate_reg_1[1146]),.o(intermediate_reg_2[573]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1145]),.i2(intermediate_reg_1[1144]),.o(intermediate_reg_2[572])); 
mux_module mux_module_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1143]),.i2(intermediate_reg_1[1142]),.o(intermediate_reg_2[571]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1141]),.i2(intermediate_reg_1[1140]),.o(intermediate_reg_2[570])); 
xor_module xor_module_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1139]),.i2(intermediate_reg_1[1138]),.o(intermediate_reg_2[569])); 
mux_module mux_module_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1137]),.i2(intermediate_reg_1[1136]),.o(intermediate_reg_2[568]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1135]),.i2(intermediate_reg_1[1134]),.o(intermediate_reg_2[567]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1133]),.i2(intermediate_reg_1[1132]),.o(intermediate_reg_2[566]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1131]),.i2(intermediate_reg_1[1130]),.o(intermediate_reg_2[565]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1129]),.i2(intermediate_reg_1[1128]),.o(intermediate_reg_2[564])); 
mux_module mux_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1127]),.i2(intermediate_reg_1[1126]),.o(intermediate_reg_2[563]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1125]),.i2(intermediate_reg_1[1124]),.o(intermediate_reg_2[562])); 
mux_module mux_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1123]),.i2(intermediate_reg_1[1122]),.o(intermediate_reg_2[561]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1121]),.i2(intermediate_reg_1[1120]),.o(intermediate_reg_2[560]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1119]),.i2(intermediate_reg_1[1118]),.o(intermediate_reg_2[559])); 
xor_module xor_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1117]),.i2(intermediate_reg_1[1116]),.o(intermediate_reg_2[558])); 
mux_module mux_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1115]),.i2(intermediate_reg_1[1114]),.o(intermediate_reg_2[557]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1113]),.i2(intermediate_reg_1[1112]),.o(intermediate_reg_2[556]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1111]),.i2(intermediate_reg_1[1110]),.o(intermediate_reg_2[555])); 
xor_module xor_module_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1109]),.i2(intermediate_reg_1[1108]),.o(intermediate_reg_2[554])); 
mux_module mux_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1107]),.i2(intermediate_reg_1[1106]),.o(intermediate_reg_2[553]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1105]),.i2(intermediate_reg_1[1104]),.o(intermediate_reg_2[552]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1103]),.i2(intermediate_reg_1[1102]),.o(intermediate_reg_2[551])); 
mux_module mux_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1101]),.i2(intermediate_reg_1[1100]),.o(intermediate_reg_2[550]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1099]),.i2(intermediate_reg_1[1098]),.o(intermediate_reg_2[549]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1097]),.i2(intermediate_reg_1[1096]),.o(intermediate_reg_2[548]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1095]),.i2(intermediate_reg_1[1094]),.o(intermediate_reg_2[547])); 
mux_module mux_module_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1093]),.i2(intermediate_reg_1[1092]),.o(intermediate_reg_2[546]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1091]),.i2(intermediate_reg_1[1090]),.o(intermediate_reg_2[545]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1089]),.i2(intermediate_reg_1[1088]),.o(intermediate_reg_2[544]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1087]),.i2(intermediate_reg_1[1086]),.o(intermediate_reg_2[543]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1085]),.i2(intermediate_reg_1[1084]),.o(intermediate_reg_2[542]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1083]),.i2(intermediate_reg_1[1082]),.o(intermediate_reg_2[541])); 
xor_module xor_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1081]),.i2(intermediate_reg_1[1080]),.o(intermediate_reg_2[540])); 
mux_module mux_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1079]),.i2(intermediate_reg_1[1078]),.o(intermediate_reg_2[539]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1077]),.i2(intermediate_reg_1[1076]),.o(intermediate_reg_2[538]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1075]),.i2(intermediate_reg_1[1074]),.o(intermediate_reg_2[537]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1073]),.i2(intermediate_reg_1[1072]),.o(intermediate_reg_2[536]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1071]),.i2(intermediate_reg_1[1070]),.o(intermediate_reg_2[535]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1069]),.i2(intermediate_reg_1[1068]),.o(intermediate_reg_2[534])); 
xor_module xor_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1067]),.i2(intermediate_reg_1[1066]),.o(intermediate_reg_2[533])); 
xor_module xor_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1065]),.i2(intermediate_reg_1[1064]),.o(intermediate_reg_2[532])); 
xor_module xor_module_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1063]),.i2(intermediate_reg_1[1062]),.o(intermediate_reg_2[531])); 
xor_module xor_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1061]),.i2(intermediate_reg_1[1060]),.o(intermediate_reg_2[530])); 
mux_module mux_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1059]),.i2(intermediate_reg_1[1058]),.o(intermediate_reg_2[529]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1057]),.i2(intermediate_reg_1[1056]),.o(intermediate_reg_2[528]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1055]),.i2(intermediate_reg_1[1054]),.o(intermediate_reg_2[527])); 
mux_module mux_module_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1053]),.i2(intermediate_reg_1[1052]),.o(intermediate_reg_2[526]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1051]),.i2(intermediate_reg_1[1050]),.o(intermediate_reg_2[525]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1049]),.i2(intermediate_reg_1[1048]),.o(intermediate_reg_2[524])); 
mux_module mux_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1047]),.i2(intermediate_reg_1[1046]),.o(intermediate_reg_2[523]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1045]),.i2(intermediate_reg_1[1044]),.o(intermediate_reg_2[522])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1043]),.i2(intermediate_reg_1[1042]),.o(intermediate_reg_2[521]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1041]),.i2(intermediate_reg_1[1040]),.o(intermediate_reg_2[520])); 
mux_module mux_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1039]),.i2(intermediate_reg_1[1038]),.o(intermediate_reg_2[519]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1037]),.i2(intermediate_reg_1[1036]),.o(intermediate_reg_2[518])); 
xor_module xor_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1035]),.i2(intermediate_reg_1[1034]),.o(intermediate_reg_2[517])); 
xor_module xor_module_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1033]),.i2(intermediate_reg_1[1032]),.o(intermediate_reg_2[516])); 
xor_module xor_module_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1031]),.i2(intermediate_reg_1[1030]),.o(intermediate_reg_2[515])); 
mux_module mux_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1029]),.i2(intermediate_reg_1[1028]),.o(intermediate_reg_2[514]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512])); 
xor_module xor_module_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511])); 
xor_module xor_module_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510])); 
mux_module mux_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508])); 
mux_module mux_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505])); 
xor_module xor_module_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504])); 
xor_module xor_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503])); 
mux_module mux_module_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501])); 
xor_module xor_module_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500])); 
mux_module mux_module_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497])); 
xor_module xor_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496])); 
xor_module xor_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495])); 
mux_module mux_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493])); 
mux_module mux_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491])); 
mux_module mux_module_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486])); 
mux_module mux_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481])); 
mux_module mux_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476])); 
xor_module xor_module_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475])); 
mux_module mux_module_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473])); 
mux_module mux_module_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470])); 
mux_module mux_module_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467])); 
mux_module mux_module_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465])); 
mux_module mux_module_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463])); 
mux_module mux_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460])); 
xor_module xor_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459])); 
xor_module xor_module_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458])); 
mux_module mux_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456])); 
xor_module xor_module_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455])); 
mux_module mux_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453])); 
xor_module xor_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452])); 
xor_module xor_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451])); 
mux_module mux_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448])); 
mux_module mux_module_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443])); 
mux_module mux_module_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440])); 
xor_module xor_module_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439])); 
mux_module mux_module_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436])); 
xor_module xor_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435])); 
mux_module mux_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433])); 
mux_module mux_module_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430])); 
xor_module xor_module_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429])); 
xor_module xor_module_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428])); 
xor_module xor_module_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427])); 
mux_module mux_module_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424])); 
xor_module xor_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423])); 
mux_module mux_module_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419])); 
mux_module mux_module_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413])); 
xor_module xor_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412])); 
mux_module mux_module_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407])); 
mux_module mux_module_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404])); 
xor_module xor_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403])); 
mux_module mux_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401])); 
xor_module xor_module_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400])); 
xor_module xor_module_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399])); 
xor_module xor_module_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398])); 
mux_module mux_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395])); 
mux_module mux_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391])); 
xor_module xor_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390])); 
xor_module xor_module_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389])); 
mux_module mux_module_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384])); 
xor_module xor_module_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383])); 
mux_module mux_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
mux_module mux_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379])); 
xor_module xor_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378])); 
xor_module xor_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377])); 
xor_module xor_module_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376])); 
mux_module mux_module_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373])); 
xor_module xor_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372])); 
mux_module mux_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368])); 
xor_module xor_module_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367])); 
mux_module mux_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
xor_module xor_module_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363])); 
xor_module xor_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362])); 
mux_module mux_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
mux_module mux_module_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357])); 
mux_module mux_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353])); 
xor_module xor_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352])); 
mux_module mux_module_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350])); 
mux_module mux_module_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348])); 
xor_module xor_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
mux_module mux_module_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345])); 
xor_module xor_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
xor_module xor_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343])); 
xor_module xor_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342])); 
xor_module xor_module_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341])); 
mux_module mux_module_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
xor_module xor_module_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334])); 
xor_module xor_module_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333])); 
mux_module mux_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331])); 
xor_module xor_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
mux_module mux_module_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
xor_module xor_module_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326])); 
xor_module xor_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325])); 
mux_module mux_module_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323])); 
xor_module xor_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322])); 
mux_module mux_module_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
xor_module xor_module_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319])); 
mux_module mux_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316])); 
xor_module xor_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315])); 
mux_module mux_module_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313])); 
xor_module xor_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312])); 
xor_module xor_module_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311])); 
mux_module mux_module_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309])); 
mux_module mux_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307])); 
mux_module mux_module_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305])); 
mux_module mux_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
mux_module mux_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
mux_module mux_module_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299])); 
mux_module mux_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297])); 
xor_module xor_module_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
xor_module xor_module_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
xor_module xor_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294])); 
xor_module xor_module_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
mux_module mux_module_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290])); 
xor_module xor_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289])); 
xor_module xor_module_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288])); 
xor_module xor_module_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287])); 
mux_module mux_module_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284])); 
xor_module xor_module_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
xor_module xor_module_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282])); 
mux_module mux_module_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279])); 
xor_module xor_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278])); 
mux_module mux_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
xor_module xor_module_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
xor_module xor_module_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
xor_module xor_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
mux_module mux_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
mux_module mux_module_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266])); 
xor_module xor_module_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
mux_module mux_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263])); 
xor_module xor_module_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
xor_module xor_module_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261])); 
xor_module xor_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
mux_module mux_module_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
mux_module mux_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254])); 
xor_module xor_module_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253])); 
mux_module mux_module_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250])); 
xor_module xor_module_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
mux_module mux_module_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246])); 
mux_module mux_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244])); 
xor_module xor_module_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243])); 
mux_module mux_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240])); 
xor_module xor_module_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239])); 
xor_module xor_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
mux_module mux_module_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236])); 
mux_module mux_module_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
xor_module xor_module_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233])); 
xor_module xor_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232])); 
xor_module xor_module_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231])); 
xor_module xor_module_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230])); 
mux_module mux_module_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227])); 
xor_module xor_module_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
mux_module mux_module_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224])); 
mux_module mux_module_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
mux_module mux_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220])); 
mux_module mux_module_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
mux_module mux_module_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216])); 
mux_module mux_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
xor_module xor_module_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
mux_module mux_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
mux_module mux_module_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
xor_module xor_module_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
xor_module xor_module_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
mux_module mux_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202])); 
xor_module xor_module_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201])); 
mux_module mux_module_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198])); 
mux_module mux_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
xor_module xor_module_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195])); 
mux_module mux_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193])); 
xor_module xor_module_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
xor_module xor_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
mux_module mux_module_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189])); 
xor_module xor_module_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
xor_module xor_module_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
mux_module mux_module_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185])); 
mux_module mux_module_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178])); 
xor_module xor_module_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
mux_module mux_module_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175])); 
mux_module mux_module_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
xor_module xor_module_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
xor_module xor_module_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
xor_module xor_module_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
xor_module xor_module_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169])); 
mux_module mux_module_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167])); 
xor_module xor_module_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166])); 
xor_module xor_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
mux_module mux_module_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
mux_module mux_module_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161])); 
mux_module mux_module_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
xor_module xor_module_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158])); 
xor_module xor_module_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157])); 
xor_module xor_module_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156])); 
mux_module mux_module_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152])); 
mux_module mux_module_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
xor_module xor_module_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
mux_module mux_module_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139])); 
mux_module mux_module_inst_2_517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
xor_module xor_module_inst_2_522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133])); 
xor_module xor_module_inst_2_523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132])); 
xor_module xor_module_inst_2_524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131])); 
xor_module xor_module_inst_2_525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130])); 
mux_module mux_module_inst_2_526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
xor_module xor_module_inst_2_528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
mux_module mux_module_inst_2_529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
xor_module xor_module_inst_2_531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124])); 
mux_module mux_module_inst_2_532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
mux_module mux_module_inst_2_534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120])); 
mux_module mux_module_inst_2_536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116])); 
xor_module xor_module_inst_2_540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115])); 
xor_module xor_module_inst_2_541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
xor_module xor_module_inst_2_542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113])); 
xor_module xor_module_inst_2_543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
mux_module mux_module_inst_2_544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
xor_module xor_module_inst_2_546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
xor_module xor_module_inst_2_547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
mux_module mux_module_inst_2_548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105])); 
xor_module xor_module_inst_2_551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104])); 
mux_module mux_module_inst_2_552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
mux_module mux_module_inst_2_555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99])); 
xor_module xor_module_inst_2_557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98])); 
xor_module xor_module_inst_2_558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
xor_module xor_module_inst_2_559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96])); 
xor_module xor_module_inst_2_560(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95])); 
xor_module xor_module_inst_2_561(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94])); 
xor_module xor_module_inst_2_562(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
xor_module xor_module_inst_2_563(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92])); 
xor_module xor_module_inst_2_564(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91])); 
xor_module xor_module_inst_2_565(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
mux_module mux_module_inst_2_566(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_567(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_568(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
mux_module mux_module_inst_2_569(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_570(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
mux_module mux_module_inst_2_571(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_572(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
mux_module mux_module_inst_2_573(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_574(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
mux_module mux_module_inst_2_575(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_576(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_577(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_578(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
xor_module xor_module_inst_2_579(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76])); 
xor_module xor_module_inst_2_580(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
mux_module mux_module_inst_2_581(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_582(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73])); 
xor_module xor_module_inst_2_583(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72])); 
mux_module mux_module_inst_2_584(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_585(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_586(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_587(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68])); 
xor_module xor_module_inst_2_588(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67])); 
mux_module mux_module_inst_2_589(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_590(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65])); 
xor_module xor_module_inst_2_591(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64])); 
xor_module xor_module_inst_2_592(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
xor_module xor_module_inst_2_593(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
xor_module xor_module_inst_2_594(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
xor_module xor_module_inst_2_595(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60])); 
mux_module mux_module_inst_2_596(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_597(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
xor_module xor_module_inst_2_598(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57])); 
mux_module mux_module_inst_2_599(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_600(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_601(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54])); 
mux_module mux_module_inst_2_602(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_603(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_604(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_605(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
xor_module xor_module_inst_2_606(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
mux_module mux_module_inst_2_607(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_608(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_609(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46])); 
xor_module xor_module_inst_2_610(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45])); 
xor_module xor_module_inst_2_611(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44])); 
mux_module mux_module_inst_2_612(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_613(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_614(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_615(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_616(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39])); 
xor_module xor_module_inst_2_617(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38])); 
mux_module mux_module_inst_2_618(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_619(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_620(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_621(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_622(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_623(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_624(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_625(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_626(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_627(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
mux_module mux_module_inst_2_628(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_629(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_630(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_631(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
mux_module mux_module_inst_2_632(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_633(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_634(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_635(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_636(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
mux_module mux_module_inst_2_637(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_638(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_639(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_640(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15])); 
mux_module mux_module_inst_2_641(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_642(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13])); 
mux_module mux_module_inst_2_643(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_644(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_645(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10])); 
xor_module xor_module_inst_2_646(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
xor_module xor_module_inst_2_647(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8])); 
mux_module mux_module_inst_2_648(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_649(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_650(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_651(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_652(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
mux_module mux_module_inst_2_653(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_654(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_655(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0]),.sel(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [655:0] <= intermediate_reg_2; 
outp[1055:656] <= intermediate_reg_2[399:0] ; 
end 
endmodule 
 

module interface_12(input [303:0] inp, output reg [511:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[303:0] <= inp ; 
outp[511:304] <= inp[207:0] ; 
end 
endmodule 

module interface_13(input [4143:0] inp, output reg [1319:0] outp, input clk, input reset);
reg [4143:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [2071:0]intermediate_reg_1; 
 
xor_module xor_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4143]),.i2(intermediate_reg_0[4142]),.o(intermediate_reg_1[2071])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4141]),.i2(intermediate_reg_0[4140]),.o(intermediate_reg_1[2070]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4139]),.i2(intermediate_reg_0[4138]),.o(intermediate_reg_1[2069]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4137]),.i2(intermediate_reg_0[4136]),.o(intermediate_reg_1[2068])); 
xor_module xor_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4135]),.i2(intermediate_reg_0[4134]),.o(intermediate_reg_1[2067])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4133]),.i2(intermediate_reg_0[4132]),.o(intermediate_reg_1[2066])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4131]),.i2(intermediate_reg_0[4130]),.o(intermediate_reg_1[2065]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4129]),.i2(intermediate_reg_0[4128]),.o(intermediate_reg_1[2064]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4127]),.i2(intermediate_reg_0[4126]),.o(intermediate_reg_1[2063]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4125]),.i2(intermediate_reg_0[4124]),.o(intermediate_reg_1[2062]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4123]),.i2(intermediate_reg_0[4122]),.o(intermediate_reg_1[2061])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4121]),.i2(intermediate_reg_0[4120]),.o(intermediate_reg_1[2060]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4119]),.i2(intermediate_reg_0[4118]),.o(intermediate_reg_1[2059]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4117]),.i2(intermediate_reg_0[4116]),.o(intermediate_reg_1[2058])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4115]),.i2(intermediate_reg_0[4114]),.o(intermediate_reg_1[2057])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4113]),.i2(intermediate_reg_0[4112]),.o(intermediate_reg_1[2056]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4111]),.i2(intermediate_reg_0[4110]),.o(intermediate_reg_1[2055]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4109]),.i2(intermediate_reg_0[4108]),.o(intermediate_reg_1[2054])); 
xor_module xor_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4107]),.i2(intermediate_reg_0[4106]),.o(intermediate_reg_1[2053])); 
xor_module xor_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4105]),.i2(intermediate_reg_0[4104]),.o(intermediate_reg_1[2052])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4103]),.i2(intermediate_reg_0[4102]),.o(intermediate_reg_1[2051])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4101]),.i2(intermediate_reg_0[4100]),.o(intermediate_reg_1[2050])); 
xor_module xor_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4099]),.i2(intermediate_reg_0[4098]),.o(intermediate_reg_1[2049])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4097]),.i2(intermediate_reg_0[4096]),.o(intermediate_reg_1[2048])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4095]),.i2(intermediate_reg_0[4094]),.o(intermediate_reg_1[2047]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4093]),.i2(intermediate_reg_0[4092]),.o(intermediate_reg_1[2046]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4091]),.i2(intermediate_reg_0[4090]),.o(intermediate_reg_1[2045])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4089]),.i2(intermediate_reg_0[4088]),.o(intermediate_reg_1[2044])); 
xor_module xor_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4087]),.i2(intermediate_reg_0[4086]),.o(intermediate_reg_1[2043])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4085]),.i2(intermediate_reg_0[4084]),.o(intermediate_reg_1[2042]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4083]),.i2(intermediate_reg_0[4082]),.o(intermediate_reg_1[2041])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4081]),.i2(intermediate_reg_0[4080]),.o(intermediate_reg_1[2040]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4079]),.i2(intermediate_reg_0[4078]),.o(intermediate_reg_1[2039])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4077]),.i2(intermediate_reg_0[4076]),.o(intermediate_reg_1[2038]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4075]),.i2(intermediate_reg_0[4074]),.o(intermediate_reg_1[2037]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4073]),.i2(intermediate_reg_0[4072]),.o(intermediate_reg_1[2036])); 
xor_module xor_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4071]),.i2(intermediate_reg_0[4070]),.o(intermediate_reg_1[2035])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4069]),.i2(intermediate_reg_0[4068]),.o(intermediate_reg_1[2034])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4067]),.i2(intermediate_reg_0[4066]),.o(intermediate_reg_1[2033])); 
xor_module xor_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4065]),.i2(intermediate_reg_0[4064]),.o(intermediate_reg_1[2032])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4063]),.i2(intermediate_reg_0[4062]),.o(intermediate_reg_1[2031])); 
mux_module mux_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4061]),.i2(intermediate_reg_0[4060]),.o(intermediate_reg_1[2030]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4059]),.i2(intermediate_reg_0[4058]),.o(intermediate_reg_1[2029])); 
mux_module mux_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4057]),.i2(intermediate_reg_0[4056]),.o(intermediate_reg_1[2028]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4055]),.i2(intermediate_reg_0[4054]),.o(intermediate_reg_1[2027]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4053]),.i2(intermediate_reg_0[4052]),.o(intermediate_reg_1[2026])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4051]),.i2(intermediate_reg_0[4050]),.o(intermediate_reg_1[2025]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4049]),.i2(intermediate_reg_0[4048]),.o(intermediate_reg_1[2024]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4047]),.i2(intermediate_reg_0[4046]),.o(intermediate_reg_1[2023])); 
xor_module xor_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4045]),.i2(intermediate_reg_0[4044]),.o(intermediate_reg_1[2022])); 
xor_module xor_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4043]),.i2(intermediate_reg_0[4042]),.o(intermediate_reg_1[2021])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4041]),.i2(intermediate_reg_0[4040]),.o(intermediate_reg_1[2020])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4039]),.i2(intermediate_reg_0[4038]),.o(intermediate_reg_1[2019]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4037]),.i2(intermediate_reg_0[4036]),.o(intermediate_reg_1[2018]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4035]),.i2(intermediate_reg_0[4034]),.o(intermediate_reg_1[2017])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4033]),.i2(intermediate_reg_0[4032]),.o(intermediate_reg_1[2016]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4031]),.i2(intermediate_reg_0[4030]),.o(intermediate_reg_1[2015])); 
xor_module xor_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4029]),.i2(intermediate_reg_0[4028]),.o(intermediate_reg_1[2014])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4027]),.i2(intermediate_reg_0[4026]),.o(intermediate_reg_1[2013])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4025]),.i2(intermediate_reg_0[4024]),.o(intermediate_reg_1[2012])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4023]),.i2(intermediate_reg_0[4022]),.o(intermediate_reg_1[2011])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4021]),.i2(intermediate_reg_0[4020]),.o(intermediate_reg_1[2010])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4019]),.i2(intermediate_reg_0[4018]),.o(intermediate_reg_1[2009]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4017]),.i2(intermediate_reg_0[4016]),.o(intermediate_reg_1[2008])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4015]),.i2(intermediate_reg_0[4014]),.o(intermediate_reg_1[2007])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4013]),.i2(intermediate_reg_0[4012]),.o(intermediate_reg_1[2006])); 
xor_module xor_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4011]),.i2(intermediate_reg_0[4010]),.o(intermediate_reg_1[2005])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4009]),.i2(intermediate_reg_0[4008]),.o(intermediate_reg_1[2004])); 
xor_module xor_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4007]),.i2(intermediate_reg_0[4006]),.o(intermediate_reg_1[2003])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4005]),.i2(intermediate_reg_0[4004]),.o(intermediate_reg_1[2002])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4003]),.i2(intermediate_reg_0[4002]),.o(intermediate_reg_1[2001])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4001]),.i2(intermediate_reg_0[4000]),.o(intermediate_reg_1[2000]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3999]),.i2(intermediate_reg_0[3998]),.o(intermediate_reg_1[1999]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3997]),.i2(intermediate_reg_0[3996]),.o(intermediate_reg_1[1998])); 
xor_module xor_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3995]),.i2(intermediate_reg_0[3994]),.o(intermediate_reg_1[1997])); 
xor_module xor_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3993]),.i2(intermediate_reg_0[3992]),.o(intermediate_reg_1[1996])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3991]),.i2(intermediate_reg_0[3990]),.o(intermediate_reg_1[1995])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3989]),.i2(intermediate_reg_0[3988]),.o(intermediate_reg_1[1994]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3987]),.i2(intermediate_reg_0[3986]),.o(intermediate_reg_1[1993]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3985]),.i2(intermediate_reg_0[3984]),.o(intermediate_reg_1[1992])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3983]),.i2(intermediate_reg_0[3982]),.o(intermediate_reg_1[1991])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3981]),.i2(intermediate_reg_0[3980]),.o(intermediate_reg_1[1990])); 
xor_module xor_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3979]),.i2(intermediate_reg_0[3978]),.o(intermediate_reg_1[1989])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3977]),.i2(intermediate_reg_0[3976]),.o(intermediate_reg_1[1988])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3975]),.i2(intermediate_reg_0[3974]),.o(intermediate_reg_1[1987]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3973]),.i2(intermediate_reg_0[3972]),.o(intermediate_reg_1[1986]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3971]),.i2(intermediate_reg_0[3970]),.o(intermediate_reg_1[1985])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3969]),.i2(intermediate_reg_0[3968]),.o(intermediate_reg_1[1984])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3967]),.i2(intermediate_reg_0[3966]),.o(intermediate_reg_1[1983])); 
mux_module mux_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3965]),.i2(intermediate_reg_0[3964]),.o(intermediate_reg_1[1982]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3963]),.i2(intermediate_reg_0[3962]),.o(intermediate_reg_1[1981])); 
xor_module xor_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3961]),.i2(intermediate_reg_0[3960]),.o(intermediate_reg_1[1980])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3959]),.i2(intermediate_reg_0[3958]),.o(intermediate_reg_1[1979])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3957]),.i2(intermediate_reg_0[3956]),.o(intermediate_reg_1[1978])); 
xor_module xor_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3955]),.i2(intermediate_reg_0[3954]),.o(intermediate_reg_1[1977])); 
xor_module xor_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3953]),.i2(intermediate_reg_0[3952]),.o(intermediate_reg_1[1976])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3951]),.i2(intermediate_reg_0[3950]),.o(intermediate_reg_1[1975])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3949]),.i2(intermediate_reg_0[3948]),.o(intermediate_reg_1[1974]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3947]),.i2(intermediate_reg_0[3946]),.o(intermediate_reg_1[1973])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3945]),.i2(intermediate_reg_0[3944]),.o(intermediate_reg_1[1972])); 
xor_module xor_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3943]),.i2(intermediate_reg_0[3942]),.o(intermediate_reg_1[1971])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3941]),.i2(intermediate_reg_0[3940]),.o(intermediate_reg_1[1970])); 
xor_module xor_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3939]),.i2(intermediate_reg_0[3938]),.o(intermediate_reg_1[1969])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3937]),.i2(intermediate_reg_0[3936]),.o(intermediate_reg_1[1968]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3935]),.i2(intermediate_reg_0[3934]),.o(intermediate_reg_1[1967]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3933]),.i2(intermediate_reg_0[3932]),.o(intermediate_reg_1[1966])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3931]),.i2(intermediate_reg_0[3930]),.o(intermediate_reg_1[1965])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3929]),.i2(intermediate_reg_0[3928]),.o(intermediate_reg_1[1964]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3927]),.i2(intermediate_reg_0[3926]),.o(intermediate_reg_1[1963]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3925]),.i2(intermediate_reg_0[3924]),.o(intermediate_reg_1[1962])); 
xor_module xor_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3923]),.i2(intermediate_reg_0[3922]),.o(intermediate_reg_1[1961])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3921]),.i2(intermediate_reg_0[3920]),.o(intermediate_reg_1[1960]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3919]),.i2(intermediate_reg_0[3918]),.o(intermediate_reg_1[1959])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3917]),.i2(intermediate_reg_0[3916]),.o(intermediate_reg_1[1958])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3915]),.i2(intermediate_reg_0[3914]),.o(intermediate_reg_1[1957]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3913]),.i2(intermediate_reg_0[3912]),.o(intermediate_reg_1[1956]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3911]),.i2(intermediate_reg_0[3910]),.o(intermediate_reg_1[1955]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3909]),.i2(intermediate_reg_0[3908]),.o(intermediate_reg_1[1954])); 
xor_module xor_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3907]),.i2(intermediate_reg_0[3906]),.o(intermediate_reg_1[1953])); 
xor_module xor_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3905]),.i2(intermediate_reg_0[3904]),.o(intermediate_reg_1[1952])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3903]),.i2(intermediate_reg_0[3902]),.o(intermediate_reg_1[1951]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3901]),.i2(intermediate_reg_0[3900]),.o(intermediate_reg_1[1950])); 
xor_module xor_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3899]),.i2(intermediate_reg_0[3898]),.o(intermediate_reg_1[1949])); 
xor_module xor_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3897]),.i2(intermediate_reg_0[3896]),.o(intermediate_reg_1[1948])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3895]),.i2(intermediate_reg_0[3894]),.o(intermediate_reg_1[1947]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3893]),.i2(intermediate_reg_0[3892]),.o(intermediate_reg_1[1946]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3891]),.i2(intermediate_reg_0[3890]),.o(intermediate_reg_1[1945])); 
xor_module xor_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3889]),.i2(intermediate_reg_0[3888]),.o(intermediate_reg_1[1944])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3887]),.i2(intermediate_reg_0[3886]),.o(intermediate_reg_1[1943]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3885]),.i2(intermediate_reg_0[3884]),.o(intermediate_reg_1[1942])); 
xor_module xor_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3883]),.i2(intermediate_reg_0[3882]),.o(intermediate_reg_1[1941])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3881]),.i2(intermediate_reg_0[3880]),.o(intermediate_reg_1[1940])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3879]),.i2(intermediate_reg_0[3878]),.o(intermediate_reg_1[1939]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3877]),.i2(intermediate_reg_0[3876]),.o(intermediate_reg_1[1938])); 
xor_module xor_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3875]),.i2(intermediate_reg_0[3874]),.o(intermediate_reg_1[1937])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3873]),.i2(intermediate_reg_0[3872]),.o(intermediate_reg_1[1936]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3871]),.i2(intermediate_reg_0[3870]),.o(intermediate_reg_1[1935])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3869]),.i2(intermediate_reg_0[3868]),.o(intermediate_reg_1[1934])); 
xor_module xor_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3867]),.i2(intermediate_reg_0[3866]),.o(intermediate_reg_1[1933])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3865]),.i2(intermediate_reg_0[3864]),.o(intermediate_reg_1[1932])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3863]),.i2(intermediate_reg_0[3862]),.o(intermediate_reg_1[1931])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3861]),.i2(intermediate_reg_0[3860]),.o(intermediate_reg_1[1930])); 
mux_module mux_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3859]),.i2(intermediate_reg_0[3858]),.o(intermediate_reg_1[1929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3857]),.i2(intermediate_reg_0[3856]),.o(intermediate_reg_1[1928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3855]),.i2(intermediate_reg_0[3854]),.o(intermediate_reg_1[1927]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3853]),.i2(intermediate_reg_0[3852]),.o(intermediate_reg_1[1926])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3851]),.i2(intermediate_reg_0[3850]),.o(intermediate_reg_1[1925]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3849]),.i2(intermediate_reg_0[3848]),.o(intermediate_reg_1[1924])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3847]),.i2(intermediate_reg_0[3846]),.o(intermediate_reg_1[1923]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3845]),.i2(intermediate_reg_0[3844]),.o(intermediate_reg_1[1922])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3843]),.i2(intermediate_reg_0[3842]),.o(intermediate_reg_1[1921]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3841]),.i2(intermediate_reg_0[3840]),.o(intermediate_reg_1[1920])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3839]),.i2(intermediate_reg_0[3838]),.o(intermediate_reg_1[1919])); 
xor_module xor_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3837]),.i2(intermediate_reg_0[3836]),.o(intermediate_reg_1[1918])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3835]),.i2(intermediate_reg_0[3834]),.o(intermediate_reg_1[1917]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3833]),.i2(intermediate_reg_0[3832]),.o(intermediate_reg_1[1916])); 
xor_module xor_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3831]),.i2(intermediate_reg_0[3830]),.o(intermediate_reg_1[1915])); 
mux_module mux_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3829]),.i2(intermediate_reg_0[3828]),.o(intermediate_reg_1[1914]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3827]),.i2(intermediate_reg_0[3826]),.o(intermediate_reg_1[1913])); 
mux_module mux_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3825]),.i2(intermediate_reg_0[3824]),.o(intermediate_reg_1[1912]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3823]),.i2(intermediate_reg_0[3822]),.o(intermediate_reg_1[1911])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3821]),.i2(intermediate_reg_0[3820]),.o(intermediate_reg_1[1910]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3819]),.i2(intermediate_reg_0[3818]),.o(intermediate_reg_1[1909])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3817]),.i2(intermediate_reg_0[3816]),.o(intermediate_reg_1[1908]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3815]),.i2(intermediate_reg_0[3814]),.o(intermediate_reg_1[1907]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3813]),.i2(intermediate_reg_0[3812]),.o(intermediate_reg_1[1906])); 
xor_module xor_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3811]),.i2(intermediate_reg_0[3810]),.o(intermediate_reg_1[1905])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3809]),.i2(intermediate_reg_0[3808]),.o(intermediate_reg_1[1904]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3807]),.i2(intermediate_reg_0[3806]),.o(intermediate_reg_1[1903])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3805]),.i2(intermediate_reg_0[3804]),.o(intermediate_reg_1[1902]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3803]),.i2(intermediate_reg_0[3802]),.o(intermediate_reg_1[1901]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3801]),.i2(intermediate_reg_0[3800]),.o(intermediate_reg_1[1900])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3799]),.i2(intermediate_reg_0[3798]),.o(intermediate_reg_1[1899])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3797]),.i2(intermediate_reg_0[3796]),.o(intermediate_reg_1[1898]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3795]),.i2(intermediate_reg_0[3794]),.o(intermediate_reg_1[1897])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3793]),.i2(intermediate_reg_0[3792]),.o(intermediate_reg_1[1896]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3791]),.i2(intermediate_reg_0[3790]),.o(intermediate_reg_1[1895])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3789]),.i2(intermediate_reg_0[3788]),.o(intermediate_reg_1[1894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3787]),.i2(intermediate_reg_0[3786]),.o(intermediate_reg_1[1893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3785]),.i2(intermediate_reg_0[3784]),.o(intermediate_reg_1[1892]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3783]),.i2(intermediate_reg_0[3782]),.o(intermediate_reg_1[1891])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3781]),.i2(intermediate_reg_0[3780]),.o(intermediate_reg_1[1890]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3779]),.i2(intermediate_reg_0[3778]),.o(intermediate_reg_1[1889])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3777]),.i2(intermediate_reg_0[3776]),.o(intermediate_reg_1[1888]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3775]),.i2(intermediate_reg_0[3774]),.o(intermediate_reg_1[1887]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3773]),.i2(intermediate_reg_0[3772]),.o(intermediate_reg_1[1886])); 
xor_module xor_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3771]),.i2(intermediate_reg_0[3770]),.o(intermediate_reg_1[1885])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3769]),.i2(intermediate_reg_0[3768]),.o(intermediate_reg_1[1884]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3767]),.i2(intermediate_reg_0[3766]),.o(intermediate_reg_1[1883])); 
xor_module xor_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3765]),.i2(intermediate_reg_0[3764]),.o(intermediate_reg_1[1882])); 
xor_module xor_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3763]),.i2(intermediate_reg_0[3762]),.o(intermediate_reg_1[1881])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3761]),.i2(intermediate_reg_0[3760]),.o(intermediate_reg_1[1880])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3759]),.i2(intermediate_reg_0[3758]),.o(intermediate_reg_1[1879])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3757]),.i2(intermediate_reg_0[3756]),.o(intermediate_reg_1[1878]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3755]),.i2(intermediate_reg_0[3754]),.o(intermediate_reg_1[1877])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3753]),.i2(intermediate_reg_0[3752]),.o(intermediate_reg_1[1876])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3751]),.i2(intermediate_reg_0[3750]),.o(intermediate_reg_1[1875]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3749]),.i2(intermediate_reg_0[3748]),.o(intermediate_reg_1[1874])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3747]),.i2(intermediate_reg_0[3746]),.o(intermediate_reg_1[1873]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3745]),.i2(intermediate_reg_0[3744]),.o(intermediate_reg_1[1872]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3743]),.i2(intermediate_reg_0[3742]),.o(intermediate_reg_1[1871])); 
xor_module xor_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3741]),.i2(intermediate_reg_0[3740]),.o(intermediate_reg_1[1870])); 
mux_module mux_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3739]),.i2(intermediate_reg_0[3738]),.o(intermediate_reg_1[1869]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3737]),.i2(intermediate_reg_0[3736]),.o(intermediate_reg_1[1868]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3735]),.i2(intermediate_reg_0[3734]),.o(intermediate_reg_1[1867]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3733]),.i2(intermediate_reg_0[3732]),.o(intermediate_reg_1[1866])); 
xor_module xor_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3731]),.i2(intermediate_reg_0[3730]),.o(intermediate_reg_1[1865])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3729]),.i2(intermediate_reg_0[3728]),.o(intermediate_reg_1[1864])); 
xor_module xor_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3727]),.i2(intermediate_reg_0[3726]),.o(intermediate_reg_1[1863])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3725]),.i2(intermediate_reg_0[3724]),.o(intermediate_reg_1[1862]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3723]),.i2(intermediate_reg_0[3722]),.o(intermediate_reg_1[1861])); 
mux_module mux_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3721]),.i2(intermediate_reg_0[3720]),.o(intermediate_reg_1[1860]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3719]),.i2(intermediate_reg_0[3718]),.o(intermediate_reg_1[1859])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3717]),.i2(intermediate_reg_0[3716]),.o(intermediate_reg_1[1858]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3715]),.i2(intermediate_reg_0[3714]),.o(intermediate_reg_1[1857]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3713]),.i2(intermediate_reg_0[3712]),.o(intermediate_reg_1[1856])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3711]),.i2(intermediate_reg_0[3710]),.o(intermediate_reg_1[1855])); 
mux_module mux_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3709]),.i2(intermediate_reg_0[3708]),.o(intermediate_reg_1[1854]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3707]),.i2(intermediate_reg_0[3706]),.o(intermediate_reg_1[1853])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3705]),.i2(intermediate_reg_0[3704]),.o(intermediate_reg_1[1852]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3703]),.i2(intermediate_reg_0[3702]),.o(intermediate_reg_1[1851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3701]),.i2(intermediate_reg_0[3700]),.o(intermediate_reg_1[1850]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3699]),.i2(intermediate_reg_0[3698]),.o(intermediate_reg_1[1849])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3697]),.i2(intermediate_reg_0[3696]),.o(intermediate_reg_1[1848])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3695]),.i2(intermediate_reg_0[3694]),.o(intermediate_reg_1[1847])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3693]),.i2(intermediate_reg_0[3692]),.o(intermediate_reg_1[1846])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3691]),.i2(intermediate_reg_0[3690]),.o(intermediate_reg_1[1845])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3689]),.i2(intermediate_reg_0[3688]),.o(intermediate_reg_1[1844])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3687]),.i2(intermediate_reg_0[3686]),.o(intermediate_reg_1[1843])); 
xor_module xor_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3685]),.i2(intermediate_reg_0[3684]),.o(intermediate_reg_1[1842])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3683]),.i2(intermediate_reg_0[3682]),.o(intermediate_reg_1[1841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3681]),.i2(intermediate_reg_0[3680]),.o(intermediate_reg_1[1840]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3679]),.i2(intermediate_reg_0[3678]),.o(intermediate_reg_1[1839])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3677]),.i2(intermediate_reg_0[3676]),.o(intermediate_reg_1[1838]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3675]),.i2(intermediate_reg_0[3674]),.o(intermediate_reg_1[1837]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3673]),.i2(intermediate_reg_0[3672]),.o(intermediate_reg_1[1836]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3671]),.i2(intermediate_reg_0[3670]),.o(intermediate_reg_1[1835])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3669]),.i2(intermediate_reg_0[3668]),.o(intermediate_reg_1[1834])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3667]),.i2(intermediate_reg_0[3666]),.o(intermediate_reg_1[1833]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3665]),.i2(intermediate_reg_0[3664]),.o(intermediate_reg_1[1832]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3663]),.i2(intermediate_reg_0[3662]),.o(intermediate_reg_1[1831])); 
xor_module xor_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3661]),.i2(intermediate_reg_0[3660]),.o(intermediate_reg_1[1830])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3659]),.i2(intermediate_reg_0[3658]),.o(intermediate_reg_1[1829]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3657]),.i2(intermediate_reg_0[3656]),.o(intermediate_reg_1[1828])); 
xor_module xor_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3655]),.i2(intermediate_reg_0[3654]),.o(intermediate_reg_1[1827])); 
mux_module mux_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3653]),.i2(intermediate_reg_0[3652]),.o(intermediate_reg_1[1826]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3651]),.i2(intermediate_reg_0[3650]),.o(intermediate_reg_1[1825]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3649]),.i2(intermediate_reg_0[3648]),.o(intermediate_reg_1[1824])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3647]),.i2(intermediate_reg_0[3646]),.o(intermediate_reg_1[1823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3645]),.i2(intermediate_reg_0[3644]),.o(intermediate_reg_1[1822]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3643]),.i2(intermediate_reg_0[3642]),.o(intermediate_reg_1[1821])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3641]),.i2(intermediate_reg_0[3640]),.o(intermediate_reg_1[1820])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3639]),.i2(intermediate_reg_0[3638]),.o(intermediate_reg_1[1819]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3637]),.i2(intermediate_reg_0[3636]),.o(intermediate_reg_1[1818]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3635]),.i2(intermediate_reg_0[3634]),.o(intermediate_reg_1[1817])); 
xor_module xor_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3633]),.i2(intermediate_reg_0[3632]),.o(intermediate_reg_1[1816])); 
xor_module xor_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3631]),.i2(intermediate_reg_0[3630]),.o(intermediate_reg_1[1815])); 
xor_module xor_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3629]),.i2(intermediate_reg_0[3628]),.o(intermediate_reg_1[1814])); 
mux_module mux_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3627]),.i2(intermediate_reg_0[3626]),.o(intermediate_reg_1[1813]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3625]),.i2(intermediate_reg_0[3624]),.o(intermediate_reg_1[1812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3623]),.i2(intermediate_reg_0[3622]),.o(intermediate_reg_1[1811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3621]),.i2(intermediate_reg_0[3620]),.o(intermediate_reg_1[1810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3619]),.i2(intermediate_reg_0[3618]),.o(intermediate_reg_1[1809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3617]),.i2(intermediate_reg_0[3616]),.o(intermediate_reg_1[1808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3615]),.i2(intermediate_reg_0[3614]),.o(intermediate_reg_1[1807]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3613]),.i2(intermediate_reg_0[3612]),.o(intermediate_reg_1[1806])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3611]),.i2(intermediate_reg_0[3610]),.o(intermediate_reg_1[1805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3609]),.i2(intermediate_reg_0[3608]),.o(intermediate_reg_1[1804]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3607]),.i2(intermediate_reg_0[3606]),.o(intermediate_reg_1[1803])); 
mux_module mux_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3605]),.i2(intermediate_reg_0[3604]),.o(intermediate_reg_1[1802]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3603]),.i2(intermediate_reg_0[3602]),.o(intermediate_reg_1[1801])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3601]),.i2(intermediate_reg_0[3600]),.o(intermediate_reg_1[1800]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3599]),.i2(intermediate_reg_0[3598]),.o(intermediate_reg_1[1799]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3597]),.i2(intermediate_reg_0[3596]),.o(intermediate_reg_1[1798])); 
xor_module xor_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3595]),.i2(intermediate_reg_0[3594]),.o(intermediate_reg_1[1797])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3593]),.i2(intermediate_reg_0[3592]),.o(intermediate_reg_1[1796]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3591]),.i2(intermediate_reg_0[3590]),.o(intermediate_reg_1[1795])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3589]),.i2(intermediate_reg_0[3588]),.o(intermediate_reg_1[1794])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3587]),.i2(intermediate_reg_0[3586]),.o(intermediate_reg_1[1793]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3585]),.i2(intermediate_reg_0[3584]),.o(intermediate_reg_1[1792])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3583]),.i2(intermediate_reg_0[3582]),.o(intermediate_reg_1[1791])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3581]),.i2(intermediate_reg_0[3580]),.o(intermediate_reg_1[1790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3579]),.i2(intermediate_reg_0[3578]),.o(intermediate_reg_1[1789]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3577]),.i2(intermediate_reg_0[3576]),.o(intermediate_reg_1[1788])); 
xor_module xor_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3575]),.i2(intermediate_reg_0[3574]),.o(intermediate_reg_1[1787])); 
xor_module xor_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3573]),.i2(intermediate_reg_0[3572]),.o(intermediate_reg_1[1786])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3571]),.i2(intermediate_reg_0[3570]),.o(intermediate_reg_1[1785])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3569]),.i2(intermediate_reg_0[3568]),.o(intermediate_reg_1[1784]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3567]),.i2(intermediate_reg_0[3566]),.o(intermediate_reg_1[1783])); 
xor_module xor_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3565]),.i2(intermediate_reg_0[3564]),.o(intermediate_reg_1[1782])); 
mux_module mux_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3563]),.i2(intermediate_reg_0[3562]),.o(intermediate_reg_1[1781]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3561]),.i2(intermediate_reg_0[3560]),.o(intermediate_reg_1[1780])); 
xor_module xor_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3559]),.i2(intermediate_reg_0[3558]),.o(intermediate_reg_1[1779])); 
xor_module xor_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3557]),.i2(intermediate_reg_0[3556]),.o(intermediate_reg_1[1778])); 
xor_module xor_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3555]),.i2(intermediate_reg_0[3554]),.o(intermediate_reg_1[1777])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3553]),.i2(intermediate_reg_0[3552]),.o(intermediate_reg_1[1776])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3551]),.i2(intermediate_reg_0[3550]),.o(intermediate_reg_1[1775])); 
mux_module mux_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3549]),.i2(intermediate_reg_0[3548]),.o(intermediate_reg_1[1774]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3547]),.i2(intermediate_reg_0[3546]),.o(intermediate_reg_1[1773])); 
mux_module mux_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3545]),.i2(intermediate_reg_0[3544]),.o(intermediate_reg_1[1772]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3543]),.i2(intermediate_reg_0[3542]),.o(intermediate_reg_1[1771]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3541]),.i2(intermediate_reg_0[3540]),.o(intermediate_reg_1[1770]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3539]),.i2(intermediate_reg_0[3538]),.o(intermediate_reg_1[1769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3537]),.i2(intermediate_reg_0[3536]),.o(intermediate_reg_1[1768]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3535]),.i2(intermediate_reg_0[3534]),.o(intermediate_reg_1[1767])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3533]),.i2(intermediate_reg_0[3532]),.o(intermediate_reg_1[1766])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3531]),.i2(intermediate_reg_0[3530]),.o(intermediate_reg_1[1765])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3529]),.i2(intermediate_reg_0[3528]),.o(intermediate_reg_1[1764]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3527]),.i2(intermediate_reg_0[3526]),.o(intermediate_reg_1[1763])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3525]),.i2(intermediate_reg_0[3524]),.o(intermediate_reg_1[1762])); 
mux_module mux_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3523]),.i2(intermediate_reg_0[3522]),.o(intermediate_reg_1[1761]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3521]),.i2(intermediate_reg_0[3520]),.o(intermediate_reg_1[1760])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3519]),.i2(intermediate_reg_0[3518]),.o(intermediate_reg_1[1759])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3517]),.i2(intermediate_reg_0[3516]),.o(intermediate_reg_1[1758])); 
xor_module xor_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3515]),.i2(intermediate_reg_0[3514]),.o(intermediate_reg_1[1757])); 
mux_module mux_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3513]),.i2(intermediate_reg_0[3512]),.o(intermediate_reg_1[1756]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3511]),.i2(intermediate_reg_0[3510]),.o(intermediate_reg_1[1755])); 
xor_module xor_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3509]),.i2(intermediate_reg_0[3508]),.o(intermediate_reg_1[1754])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3507]),.i2(intermediate_reg_0[3506]),.o(intermediate_reg_1[1753])); 
mux_module mux_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3505]),.i2(intermediate_reg_0[3504]),.o(intermediate_reg_1[1752]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3503]),.i2(intermediate_reg_0[3502]),.o(intermediate_reg_1[1751]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3501]),.i2(intermediate_reg_0[3500]),.o(intermediate_reg_1[1750])); 
xor_module xor_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3499]),.i2(intermediate_reg_0[3498]),.o(intermediate_reg_1[1749])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3497]),.i2(intermediate_reg_0[3496]),.o(intermediate_reg_1[1748]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3495]),.i2(intermediate_reg_0[3494]),.o(intermediate_reg_1[1747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3493]),.i2(intermediate_reg_0[3492]),.o(intermediate_reg_1[1746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3491]),.i2(intermediate_reg_0[3490]),.o(intermediate_reg_1[1745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3489]),.i2(intermediate_reg_0[3488]),.o(intermediate_reg_1[1744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3487]),.i2(intermediate_reg_0[3486]),.o(intermediate_reg_1[1743]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3485]),.i2(intermediate_reg_0[3484]),.o(intermediate_reg_1[1742])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3483]),.i2(intermediate_reg_0[3482]),.o(intermediate_reg_1[1741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3481]),.i2(intermediate_reg_0[3480]),.o(intermediate_reg_1[1740]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3479]),.i2(intermediate_reg_0[3478]),.o(intermediate_reg_1[1739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3477]),.i2(intermediate_reg_0[3476]),.o(intermediate_reg_1[1738]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3475]),.i2(intermediate_reg_0[3474]),.o(intermediate_reg_1[1737]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3473]),.i2(intermediate_reg_0[3472]),.o(intermediate_reg_1[1736]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3471]),.i2(intermediate_reg_0[3470]),.o(intermediate_reg_1[1735])); 
mux_module mux_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3469]),.i2(intermediate_reg_0[3468]),.o(intermediate_reg_1[1734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3467]),.i2(intermediate_reg_0[3466]),.o(intermediate_reg_1[1733]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3465]),.i2(intermediate_reg_0[3464]),.o(intermediate_reg_1[1732]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3463]),.i2(intermediate_reg_0[3462]),.o(intermediate_reg_1[1731])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3461]),.i2(intermediate_reg_0[3460]),.o(intermediate_reg_1[1730])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3459]),.i2(intermediate_reg_0[3458]),.o(intermediate_reg_1[1729]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3457]),.i2(intermediate_reg_0[3456]),.o(intermediate_reg_1[1728])); 
mux_module mux_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3455]),.i2(intermediate_reg_0[3454]),.o(intermediate_reg_1[1727]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3453]),.i2(intermediate_reg_0[3452]),.o(intermediate_reg_1[1726])); 
mux_module mux_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3451]),.i2(intermediate_reg_0[3450]),.o(intermediate_reg_1[1725]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3449]),.i2(intermediate_reg_0[3448]),.o(intermediate_reg_1[1724])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3447]),.i2(intermediate_reg_0[3446]),.o(intermediate_reg_1[1723]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3445]),.i2(intermediate_reg_0[3444]),.o(intermediate_reg_1[1722]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3443]),.i2(intermediate_reg_0[3442]),.o(intermediate_reg_1[1721])); 
mux_module mux_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3441]),.i2(intermediate_reg_0[3440]),.o(intermediate_reg_1[1720]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3439]),.i2(intermediate_reg_0[3438]),.o(intermediate_reg_1[1719]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3437]),.i2(intermediate_reg_0[3436]),.o(intermediate_reg_1[1718])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3435]),.i2(intermediate_reg_0[3434]),.o(intermediate_reg_1[1717])); 
mux_module mux_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3433]),.i2(intermediate_reg_0[3432]),.o(intermediate_reg_1[1716]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3431]),.i2(intermediate_reg_0[3430]),.o(intermediate_reg_1[1715])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3429]),.i2(intermediate_reg_0[3428]),.o(intermediate_reg_1[1714]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3427]),.i2(intermediate_reg_0[3426]),.o(intermediate_reg_1[1713]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3425]),.i2(intermediate_reg_0[3424]),.o(intermediate_reg_1[1712])); 
xor_module xor_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3423]),.i2(intermediate_reg_0[3422]),.o(intermediate_reg_1[1711])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3421]),.i2(intermediate_reg_0[3420]),.o(intermediate_reg_1[1710])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3419]),.i2(intermediate_reg_0[3418]),.o(intermediate_reg_1[1709])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3417]),.i2(intermediate_reg_0[3416]),.o(intermediate_reg_1[1708])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3415]),.i2(intermediate_reg_0[3414]),.o(intermediate_reg_1[1707])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3413]),.i2(intermediate_reg_0[3412]),.o(intermediate_reg_1[1706]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3411]),.i2(intermediate_reg_0[3410]),.o(intermediate_reg_1[1705]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3409]),.i2(intermediate_reg_0[3408]),.o(intermediate_reg_1[1704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3407]),.i2(intermediate_reg_0[3406]),.o(intermediate_reg_1[1703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3405]),.i2(intermediate_reg_0[3404]),.o(intermediate_reg_1[1702]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3403]),.i2(intermediate_reg_0[3402]),.o(intermediate_reg_1[1701])); 
xor_module xor_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3401]),.i2(intermediate_reg_0[3400]),.o(intermediate_reg_1[1700])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3399]),.i2(intermediate_reg_0[3398]),.o(intermediate_reg_1[1699])); 
xor_module xor_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3397]),.i2(intermediate_reg_0[3396]),.o(intermediate_reg_1[1698])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3395]),.i2(intermediate_reg_0[3394]),.o(intermediate_reg_1[1697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3393]),.i2(intermediate_reg_0[3392]),.o(intermediate_reg_1[1696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3391]),.i2(intermediate_reg_0[3390]),.o(intermediate_reg_1[1695])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3389]),.i2(intermediate_reg_0[3388]),.o(intermediate_reg_1[1694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3387]),.i2(intermediate_reg_0[3386]),.o(intermediate_reg_1[1693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3385]),.i2(intermediate_reg_0[3384]),.o(intermediate_reg_1[1692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3383]),.i2(intermediate_reg_0[3382]),.o(intermediate_reg_1[1691]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3381]),.i2(intermediate_reg_0[3380]),.o(intermediate_reg_1[1690])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3379]),.i2(intermediate_reg_0[3378]),.o(intermediate_reg_1[1689])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3377]),.i2(intermediate_reg_0[3376]),.o(intermediate_reg_1[1688]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3375]),.i2(intermediate_reg_0[3374]),.o(intermediate_reg_1[1687])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3373]),.i2(intermediate_reg_0[3372]),.o(intermediate_reg_1[1686]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3371]),.i2(intermediate_reg_0[3370]),.o(intermediate_reg_1[1685])); 
xor_module xor_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3369]),.i2(intermediate_reg_0[3368]),.o(intermediate_reg_1[1684])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3367]),.i2(intermediate_reg_0[3366]),.o(intermediate_reg_1[1683])); 
xor_module xor_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3365]),.i2(intermediate_reg_0[3364]),.o(intermediate_reg_1[1682])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3363]),.i2(intermediate_reg_0[3362]),.o(intermediate_reg_1[1681]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3361]),.i2(intermediate_reg_0[3360]),.o(intermediate_reg_1[1680])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3359]),.i2(intermediate_reg_0[3358]),.o(intermediate_reg_1[1679])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3357]),.i2(intermediate_reg_0[3356]),.o(intermediate_reg_1[1678]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3355]),.i2(intermediate_reg_0[3354]),.o(intermediate_reg_1[1677]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3353]),.i2(intermediate_reg_0[3352]),.o(intermediate_reg_1[1676])); 
xor_module xor_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3351]),.i2(intermediate_reg_0[3350]),.o(intermediate_reg_1[1675])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3349]),.i2(intermediate_reg_0[3348]),.o(intermediate_reg_1[1674])); 
mux_module mux_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3347]),.i2(intermediate_reg_0[3346]),.o(intermediate_reg_1[1673]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3345]),.i2(intermediate_reg_0[3344]),.o(intermediate_reg_1[1672])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3343]),.i2(intermediate_reg_0[3342]),.o(intermediate_reg_1[1671]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3341]),.i2(intermediate_reg_0[3340]),.o(intermediate_reg_1[1670])); 
mux_module mux_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3339]),.i2(intermediate_reg_0[3338]),.o(intermediate_reg_1[1669]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3337]),.i2(intermediate_reg_0[3336]),.o(intermediate_reg_1[1668])); 
mux_module mux_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3335]),.i2(intermediate_reg_0[3334]),.o(intermediate_reg_1[1667]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3333]),.i2(intermediate_reg_0[3332]),.o(intermediate_reg_1[1666])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3331]),.i2(intermediate_reg_0[3330]),.o(intermediate_reg_1[1665])); 
xor_module xor_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3329]),.i2(intermediate_reg_0[3328]),.o(intermediate_reg_1[1664])); 
mux_module mux_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3327]),.i2(intermediate_reg_0[3326]),.o(intermediate_reg_1[1663]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3325]),.i2(intermediate_reg_0[3324]),.o(intermediate_reg_1[1662]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3323]),.i2(intermediate_reg_0[3322]),.o(intermediate_reg_1[1661])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3321]),.i2(intermediate_reg_0[3320]),.o(intermediate_reg_1[1660])); 
mux_module mux_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3319]),.i2(intermediate_reg_0[3318]),.o(intermediate_reg_1[1659]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3317]),.i2(intermediate_reg_0[3316]),.o(intermediate_reg_1[1658]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3315]),.i2(intermediate_reg_0[3314]),.o(intermediate_reg_1[1657]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3313]),.i2(intermediate_reg_0[3312]),.o(intermediate_reg_1[1656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3311]),.i2(intermediate_reg_0[3310]),.o(intermediate_reg_1[1655]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3309]),.i2(intermediate_reg_0[3308]),.o(intermediate_reg_1[1654]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3307]),.i2(intermediate_reg_0[3306]),.o(intermediate_reg_1[1653]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3305]),.i2(intermediate_reg_0[3304]),.o(intermediate_reg_1[1652]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3303]),.i2(intermediate_reg_0[3302]),.o(intermediate_reg_1[1651])); 
xor_module xor_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3301]),.i2(intermediate_reg_0[3300]),.o(intermediate_reg_1[1650])); 
mux_module mux_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3299]),.i2(intermediate_reg_0[3298]),.o(intermediate_reg_1[1649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3297]),.i2(intermediate_reg_0[3296]),.o(intermediate_reg_1[1648]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3295]),.i2(intermediate_reg_0[3294]),.o(intermediate_reg_1[1647])); 
mux_module mux_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3293]),.i2(intermediate_reg_0[3292]),.o(intermediate_reg_1[1646]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3291]),.i2(intermediate_reg_0[3290]),.o(intermediate_reg_1[1645])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3289]),.i2(intermediate_reg_0[3288]),.o(intermediate_reg_1[1644]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3287]),.i2(intermediate_reg_0[3286]),.o(intermediate_reg_1[1643])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3285]),.i2(intermediate_reg_0[3284]),.o(intermediate_reg_1[1642]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3283]),.i2(intermediate_reg_0[3282]),.o(intermediate_reg_1[1641])); 
xor_module xor_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3281]),.i2(intermediate_reg_0[3280]),.o(intermediate_reg_1[1640])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3279]),.i2(intermediate_reg_0[3278]),.o(intermediate_reg_1[1639]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3277]),.i2(intermediate_reg_0[3276]),.o(intermediate_reg_1[1638])); 
xor_module xor_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3275]),.i2(intermediate_reg_0[3274]),.o(intermediate_reg_1[1637])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3273]),.i2(intermediate_reg_0[3272]),.o(intermediate_reg_1[1636])); 
xor_module xor_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3271]),.i2(intermediate_reg_0[3270]),.o(intermediate_reg_1[1635])); 
xor_module xor_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3269]),.i2(intermediate_reg_0[3268]),.o(intermediate_reg_1[1634])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3267]),.i2(intermediate_reg_0[3266]),.o(intermediate_reg_1[1633]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3265]),.i2(intermediate_reg_0[3264]),.o(intermediate_reg_1[1632])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3263]),.i2(intermediate_reg_0[3262]),.o(intermediate_reg_1[1631]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3261]),.i2(intermediate_reg_0[3260]),.o(intermediate_reg_1[1630])); 
xor_module xor_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3259]),.i2(intermediate_reg_0[3258]),.o(intermediate_reg_1[1629])); 
xor_module xor_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3257]),.i2(intermediate_reg_0[3256]),.o(intermediate_reg_1[1628])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3255]),.i2(intermediate_reg_0[3254]),.o(intermediate_reg_1[1627])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3253]),.i2(intermediate_reg_0[3252]),.o(intermediate_reg_1[1626])); 
mux_module mux_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3251]),.i2(intermediate_reg_0[3250]),.o(intermediate_reg_1[1625]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3249]),.i2(intermediate_reg_0[3248]),.o(intermediate_reg_1[1624])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3247]),.i2(intermediate_reg_0[3246]),.o(intermediate_reg_1[1623])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3245]),.i2(intermediate_reg_0[3244]),.o(intermediate_reg_1[1622]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3243]),.i2(intermediate_reg_0[3242]),.o(intermediate_reg_1[1621]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3241]),.i2(intermediate_reg_0[3240]),.o(intermediate_reg_1[1620])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3239]),.i2(intermediate_reg_0[3238]),.o(intermediate_reg_1[1619]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3237]),.i2(intermediate_reg_0[3236]),.o(intermediate_reg_1[1618])); 
xor_module xor_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3235]),.i2(intermediate_reg_0[3234]),.o(intermediate_reg_1[1617])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3233]),.i2(intermediate_reg_0[3232]),.o(intermediate_reg_1[1616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3231]),.i2(intermediate_reg_0[3230]),.o(intermediate_reg_1[1615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3229]),.i2(intermediate_reg_0[3228]),.o(intermediate_reg_1[1614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3227]),.i2(intermediate_reg_0[3226]),.o(intermediate_reg_1[1613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3225]),.i2(intermediate_reg_0[3224]),.o(intermediate_reg_1[1612]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3223]),.i2(intermediate_reg_0[3222]),.o(intermediate_reg_1[1611]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3221]),.i2(intermediate_reg_0[3220]),.o(intermediate_reg_1[1610])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3219]),.i2(intermediate_reg_0[3218]),.o(intermediate_reg_1[1609])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3217]),.i2(intermediate_reg_0[3216]),.o(intermediate_reg_1[1608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3215]),.i2(intermediate_reg_0[3214]),.o(intermediate_reg_1[1607]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3213]),.i2(intermediate_reg_0[3212]),.o(intermediate_reg_1[1606])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3211]),.i2(intermediate_reg_0[3210]),.o(intermediate_reg_1[1605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3209]),.i2(intermediate_reg_0[3208]),.o(intermediate_reg_1[1604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3207]),.i2(intermediate_reg_0[3206]),.o(intermediate_reg_1[1603]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3205]),.i2(intermediate_reg_0[3204]),.o(intermediate_reg_1[1602])); 
xor_module xor_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3203]),.i2(intermediate_reg_0[3202]),.o(intermediate_reg_1[1601])); 
xor_module xor_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3201]),.i2(intermediate_reg_0[3200]),.o(intermediate_reg_1[1600])); 
xor_module xor_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3199]),.i2(intermediate_reg_0[3198]),.o(intermediate_reg_1[1599])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3197]),.i2(intermediate_reg_0[3196]),.o(intermediate_reg_1[1598]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3195]),.i2(intermediate_reg_0[3194]),.o(intermediate_reg_1[1597])); 
xor_module xor_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3193]),.i2(intermediate_reg_0[3192]),.o(intermediate_reg_1[1596])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3191]),.i2(intermediate_reg_0[3190]),.o(intermediate_reg_1[1595]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3189]),.i2(intermediate_reg_0[3188]),.o(intermediate_reg_1[1594])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3187]),.i2(intermediate_reg_0[3186]),.o(intermediate_reg_1[1593]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3185]),.i2(intermediate_reg_0[3184]),.o(intermediate_reg_1[1592]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3183]),.i2(intermediate_reg_0[3182]),.o(intermediate_reg_1[1591]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3181]),.i2(intermediate_reg_0[3180]),.o(intermediate_reg_1[1590])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3179]),.i2(intermediate_reg_0[3178]),.o(intermediate_reg_1[1589]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3177]),.i2(intermediate_reg_0[3176]),.o(intermediate_reg_1[1588])); 
mux_module mux_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3175]),.i2(intermediate_reg_0[3174]),.o(intermediate_reg_1[1587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3173]),.i2(intermediate_reg_0[3172]),.o(intermediate_reg_1[1586]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3171]),.i2(intermediate_reg_0[3170]),.o(intermediate_reg_1[1585])); 
mux_module mux_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3169]),.i2(intermediate_reg_0[3168]),.o(intermediate_reg_1[1584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3167]),.i2(intermediate_reg_0[3166]),.o(intermediate_reg_1[1583]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3165]),.i2(intermediate_reg_0[3164]),.o(intermediate_reg_1[1582])); 
xor_module xor_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3163]),.i2(intermediate_reg_0[3162]),.o(intermediate_reg_1[1581])); 
mux_module mux_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3161]),.i2(intermediate_reg_0[3160]),.o(intermediate_reg_1[1580]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3159]),.i2(intermediate_reg_0[3158]),.o(intermediate_reg_1[1579]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3157]),.i2(intermediate_reg_0[3156]),.o(intermediate_reg_1[1578]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3155]),.i2(intermediate_reg_0[3154]),.o(intermediate_reg_1[1577])); 
mux_module mux_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3153]),.i2(intermediate_reg_0[3152]),.o(intermediate_reg_1[1576]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3151]),.i2(intermediate_reg_0[3150]),.o(intermediate_reg_1[1575])); 
xor_module xor_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3149]),.i2(intermediate_reg_0[3148]),.o(intermediate_reg_1[1574])); 
xor_module xor_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3147]),.i2(intermediate_reg_0[3146]),.o(intermediate_reg_1[1573])); 
mux_module mux_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3145]),.i2(intermediate_reg_0[3144]),.o(intermediate_reg_1[1572]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3143]),.i2(intermediate_reg_0[3142]),.o(intermediate_reg_1[1571])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3141]),.i2(intermediate_reg_0[3140]),.o(intermediate_reg_1[1570])); 
mux_module mux_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3139]),.i2(intermediate_reg_0[3138]),.o(intermediate_reg_1[1569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3137]),.i2(intermediate_reg_0[3136]),.o(intermediate_reg_1[1568]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3135]),.i2(intermediate_reg_0[3134]),.o(intermediate_reg_1[1567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3133]),.i2(intermediate_reg_0[3132]),.o(intermediate_reg_1[1566]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3131]),.i2(intermediate_reg_0[3130]),.o(intermediate_reg_1[1565])); 
xor_module xor_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3129]),.i2(intermediate_reg_0[3128]),.o(intermediate_reg_1[1564])); 
xor_module xor_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3127]),.i2(intermediate_reg_0[3126]),.o(intermediate_reg_1[1563])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3125]),.i2(intermediate_reg_0[3124]),.o(intermediate_reg_1[1562]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3123]),.i2(intermediate_reg_0[3122]),.o(intermediate_reg_1[1561]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3121]),.i2(intermediate_reg_0[3120]),.o(intermediate_reg_1[1560]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3119]),.i2(intermediate_reg_0[3118]),.o(intermediate_reg_1[1559])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3117]),.i2(intermediate_reg_0[3116]),.o(intermediate_reg_1[1558])); 
xor_module xor_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3115]),.i2(intermediate_reg_0[3114]),.o(intermediate_reg_1[1557])); 
mux_module mux_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3113]),.i2(intermediate_reg_0[3112]),.o(intermediate_reg_1[1556]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3111]),.i2(intermediate_reg_0[3110]),.o(intermediate_reg_1[1555]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3109]),.i2(intermediate_reg_0[3108]),.o(intermediate_reg_1[1554])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3107]),.i2(intermediate_reg_0[3106]),.o(intermediate_reg_1[1553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3105]),.i2(intermediate_reg_0[3104]),.o(intermediate_reg_1[1552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3103]),.i2(intermediate_reg_0[3102]),.o(intermediate_reg_1[1551]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3101]),.i2(intermediate_reg_0[3100]),.o(intermediate_reg_1[1550])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3099]),.i2(intermediate_reg_0[3098]),.o(intermediate_reg_1[1549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3097]),.i2(intermediate_reg_0[3096]),.o(intermediate_reg_1[1548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3095]),.i2(intermediate_reg_0[3094]),.o(intermediate_reg_1[1547]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3093]),.i2(intermediate_reg_0[3092]),.o(intermediate_reg_1[1546]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3091]),.i2(intermediate_reg_0[3090]),.o(intermediate_reg_1[1545])); 
mux_module mux_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3089]),.i2(intermediate_reg_0[3088]),.o(intermediate_reg_1[1544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3087]),.i2(intermediate_reg_0[3086]),.o(intermediate_reg_1[1543]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3085]),.i2(intermediate_reg_0[3084]),.o(intermediate_reg_1[1542])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3083]),.i2(intermediate_reg_0[3082]),.o(intermediate_reg_1[1541]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3081]),.i2(intermediate_reg_0[3080]),.o(intermediate_reg_1[1540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3079]),.i2(intermediate_reg_0[3078]),.o(intermediate_reg_1[1539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3077]),.i2(intermediate_reg_0[3076]),.o(intermediate_reg_1[1538]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3075]),.i2(intermediate_reg_0[3074]),.o(intermediate_reg_1[1537])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3073]),.i2(intermediate_reg_0[3072]),.o(intermediate_reg_1[1536])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3071]),.i2(intermediate_reg_0[3070]),.o(intermediate_reg_1[1535]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3069]),.i2(intermediate_reg_0[3068]),.o(intermediate_reg_1[1534]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3067]),.i2(intermediate_reg_0[3066]),.o(intermediate_reg_1[1533])); 
xor_module xor_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3065]),.i2(intermediate_reg_0[3064]),.o(intermediate_reg_1[1532])); 
xor_module xor_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3063]),.i2(intermediate_reg_0[3062]),.o(intermediate_reg_1[1531])); 
xor_module xor_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3061]),.i2(intermediate_reg_0[3060]),.o(intermediate_reg_1[1530])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3059]),.i2(intermediate_reg_0[3058]),.o(intermediate_reg_1[1529])); 
mux_module mux_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3057]),.i2(intermediate_reg_0[3056]),.o(intermediate_reg_1[1528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3055]),.i2(intermediate_reg_0[3054]),.o(intermediate_reg_1[1527]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3053]),.i2(intermediate_reg_0[3052]),.o(intermediate_reg_1[1526])); 
mux_module mux_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3051]),.i2(intermediate_reg_0[3050]),.o(intermediate_reg_1[1525]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3049]),.i2(intermediate_reg_0[3048]),.o(intermediate_reg_1[1524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3047]),.i2(intermediate_reg_0[3046]),.o(intermediate_reg_1[1523]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3045]),.i2(intermediate_reg_0[3044]),.o(intermediate_reg_1[1522])); 
xor_module xor_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3043]),.i2(intermediate_reg_0[3042]),.o(intermediate_reg_1[1521])); 
xor_module xor_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3041]),.i2(intermediate_reg_0[3040]),.o(intermediate_reg_1[1520])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3039]),.i2(intermediate_reg_0[3038]),.o(intermediate_reg_1[1519])); 
mux_module mux_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3037]),.i2(intermediate_reg_0[3036]),.o(intermediate_reg_1[1518]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3035]),.i2(intermediate_reg_0[3034]),.o(intermediate_reg_1[1517])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3033]),.i2(intermediate_reg_0[3032]),.o(intermediate_reg_1[1516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3031]),.i2(intermediate_reg_0[3030]),.o(intermediate_reg_1[1515]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3029]),.i2(intermediate_reg_0[3028]),.o(intermediate_reg_1[1514])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3027]),.i2(intermediate_reg_0[3026]),.o(intermediate_reg_1[1513])); 
mux_module mux_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3025]),.i2(intermediate_reg_0[3024]),.o(intermediate_reg_1[1512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3023]),.i2(intermediate_reg_0[3022]),.o(intermediate_reg_1[1511]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3021]),.i2(intermediate_reg_0[3020]),.o(intermediate_reg_1[1510])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3019]),.i2(intermediate_reg_0[3018]),.o(intermediate_reg_1[1509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3017]),.i2(intermediate_reg_0[3016]),.o(intermediate_reg_1[1508]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3015]),.i2(intermediate_reg_0[3014]),.o(intermediate_reg_1[1507]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3013]),.i2(intermediate_reg_0[3012]),.o(intermediate_reg_1[1506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3011]),.i2(intermediate_reg_0[3010]),.o(intermediate_reg_1[1505]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3009]),.i2(intermediate_reg_0[3008]),.o(intermediate_reg_1[1504])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3007]),.i2(intermediate_reg_0[3006]),.o(intermediate_reg_1[1503]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3005]),.i2(intermediate_reg_0[3004]),.o(intermediate_reg_1[1502])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3003]),.i2(intermediate_reg_0[3002]),.o(intermediate_reg_1[1501]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3001]),.i2(intermediate_reg_0[3000]),.o(intermediate_reg_1[1500])); 
xor_module xor_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2999]),.i2(intermediate_reg_0[2998]),.o(intermediate_reg_1[1499])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2997]),.i2(intermediate_reg_0[2996]),.o(intermediate_reg_1[1498]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2995]),.i2(intermediate_reg_0[2994]),.o(intermediate_reg_1[1497])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2993]),.i2(intermediate_reg_0[2992]),.o(intermediate_reg_1[1496]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2991]),.i2(intermediate_reg_0[2990]),.o(intermediate_reg_1[1495])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2989]),.i2(intermediate_reg_0[2988]),.o(intermediate_reg_1[1494]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2987]),.i2(intermediate_reg_0[2986]),.o(intermediate_reg_1[1493])); 
xor_module xor_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2985]),.i2(intermediate_reg_0[2984]),.o(intermediate_reg_1[1492])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2983]),.i2(intermediate_reg_0[2982]),.o(intermediate_reg_1[1491])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2981]),.i2(intermediate_reg_0[2980]),.o(intermediate_reg_1[1490])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2979]),.i2(intermediate_reg_0[2978]),.o(intermediate_reg_1[1489]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2977]),.i2(intermediate_reg_0[2976]),.o(intermediate_reg_1[1488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2975]),.i2(intermediate_reg_0[2974]),.o(intermediate_reg_1[1487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2973]),.i2(intermediate_reg_0[2972]),.o(intermediate_reg_1[1486]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2971]),.i2(intermediate_reg_0[2970]),.o(intermediate_reg_1[1485])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2969]),.i2(intermediate_reg_0[2968]),.o(intermediate_reg_1[1484])); 
xor_module xor_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2967]),.i2(intermediate_reg_0[2966]),.o(intermediate_reg_1[1483])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2965]),.i2(intermediate_reg_0[2964]),.o(intermediate_reg_1[1482])); 
mux_module mux_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2963]),.i2(intermediate_reg_0[2962]),.o(intermediate_reg_1[1481]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2961]),.i2(intermediate_reg_0[2960]),.o(intermediate_reg_1[1480])); 
xor_module xor_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2959]),.i2(intermediate_reg_0[2958]),.o(intermediate_reg_1[1479])); 
xor_module xor_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2957]),.i2(intermediate_reg_0[2956]),.o(intermediate_reg_1[1478])); 
mux_module mux_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2955]),.i2(intermediate_reg_0[2954]),.o(intermediate_reg_1[1477]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2953]),.i2(intermediate_reg_0[2952]),.o(intermediate_reg_1[1476])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2951]),.i2(intermediate_reg_0[2950]),.o(intermediate_reg_1[1475]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2949]),.i2(intermediate_reg_0[2948]),.o(intermediate_reg_1[1474])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2947]),.i2(intermediate_reg_0[2946]),.o(intermediate_reg_1[1473]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2945]),.i2(intermediate_reg_0[2944]),.o(intermediate_reg_1[1472])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2943]),.i2(intermediate_reg_0[2942]),.o(intermediate_reg_1[1471])); 
xor_module xor_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2941]),.i2(intermediate_reg_0[2940]),.o(intermediate_reg_1[1470])); 
xor_module xor_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2939]),.i2(intermediate_reg_0[2938]),.o(intermediate_reg_1[1469])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2937]),.i2(intermediate_reg_0[2936]),.o(intermediate_reg_1[1468]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2935]),.i2(intermediate_reg_0[2934]),.o(intermediate_reg_1[1467])); 
xor_module xor_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2933]),.i2(intermediate_reg_0[2932]),.o(intermediate_reg_1[1466])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2931]),.i2(intermediate_reg_0[2930]),.o(intermediate_reg_1[1465])); 
mux_module mux_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2929]),.i2(intermediate_reg_0[2928]),.o(intermediate_reg_1[1464]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2927]),.i2(intermediate_reg_0[2926]),.o(intermediate_reg_1[1463])); 
xor_module xor_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2925]),.i2(intermediate_reg_0[2924]),.o(intermediate_reg_1[1462])); 
xor_module xor_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2923]),.i2(intermediate_reg_0[2922]),.o(intermediate_reg_1[1461])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2921]),.i2(intermediate_reg_0[2920]),.o(intermediate_reg_1[1460]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2919]),.i2(intermediate_reg_0[2918]),.o(intermediate_reg_1[1459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2917]),.i2(intermediate_reg_0[2916]),.o(intermediate_reg_1[1458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2915]),.i2(intermediate_reg_0[2914]),.o(intermediate_reg_1[1457])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2913]),.i2(intermediate_reg_0[2912]),.o(intermediate_reg_1[1456]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2911]),.i2(intermediate_reg_0[2910]),.o(intermediate_reg_1[1455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2909]),.i2(intermediate_reg_0[2908]),.o(intermediate_reg_1[1454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2907]),.i2(intermediate_reg_0[2906]),.o(intermediate_reg_1[1453]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2905]),.i2(intermediate_reg_0[2904]),.o(intermediate_reg_1[1452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2903]),.i2(intermediate_reg_0[2902]),.o(intermediate_reg_1[1451]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2901]),.i2(intermediate_reg_0[2900]),.o(intermediate_reg_1[1450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2899]),.i2(intermediate_reg_0[2898]),.o(intermediate_reg_1[1449]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2897]),.i2(intermediate_reg_0[2896]),.o(intermediate_reg_1[1448]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2895]),.i2(intermediate_reg_0[2894]),.o(intermediate_reg_1[1447])); 
xor_module xor_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2893]),.i2(intermediate_reg_0[2892]),.o(intermediate_reg_1[1446])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2891]),.i2(intermediate_reg_0[2890]),.o(intermediate_reg_1[1445])); 
xor_module xor_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2889]),.i2(intermediate_reg_0[2888]),.o(intermediate_reg_1[1444])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2887]),.i2(intermediate_reg_0[2886]),.o(intermediate_reg_1[1443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2885]),.i2(intermediate_reg_0[2884]),.o(intermediate_reg_1[1442]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2883]),.i2(intermediate_reg_0[2882]),.o(intermediate_reg_1[1441]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2881]),.i2(intermediate_reg_0[2880]),.o(intermediate_reg_1[1440]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2879]),.i2(intermediate_reg_0[2878]),.o(intermediate_reg_1[1439])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2877]),.i2(intermediate_reg_0[2876]),.o(intermediate_reg_1[1438]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2875]),.i2(intermediate_reg_0[2874]),.o(intermediate_reg_1[1437])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2873]),.i2(intermediate_reg_0[2872]),.o(intermediate_reg_1[1436])); 
mux_module mux_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2871]),.i2(intermediate_reg_0[2870]),.o(intermediate_reg_1[1435]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2869]),.i2(intermediate_reg_0[2868]),.o(intermediate_reg_1[1434])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2867]),.i2(intermediate_reg_0[2866]),.o(intermediate_reg_1[1433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2865]),.i2(intermediate_reg_0[2864]),.o(intermediate_reg_1[1432]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2863]),.i2(intermediate_reg_0[2862]),.o(intermediate_reg_1[1431])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2861]),.i2(intermediate_reg_0[2860]),.o(intermediate_reg_1[1430])); 
mux_module mux_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2859]),.i2(intermediate_reg_0[2858]),.o(intermediate_reg_1[1429]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2857]),.i2(intermediate_reg_0[2856]),.o(intermediate_reg_1[1428])); 
xor_module xor_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2855]),.i2(intermediate_reg_0[2854]),.o(intermediate_reg_1[1427])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2853]),.i2(intermediate_reg_0[2852]),.o(intermediate_reg_1[1426]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2851]),.i2(intermediate_reg_0[2850]),.o(intermediate_reg_1[1425])); 
xor_module xor_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2849]),.i2(intermediate_reg_0[2848]),.o(intermediate_reg_1[1424])); 
mux_module mux_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2847]),.i2(intermediate_reg_0[2846]),.o(intermediate_reg_1[1423]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2845]),.i2(intermediate_reg_0[2844]),.o(intermediate_reg_1[1422])); 
xor_module xor_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2843]),.i2(intermediate_reg_0[2842]),.o(intermediate_reg_1[1421])); 
xor_module xor_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2841]),.i2(intermediate_reg_0[2840]),.o(intermediate_reg_1[1420])); 
mux_module mux_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2839]),.i2(intermediate_reg_0[2838]),.o(intermediate_reg_1[1419]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2837]),.i2(intermediate_reg_0[2836]),.o(intermediate_reg_1[1418])); 
xor_module xor_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2835]),.i2(intermediate_reg_0[2834]),.o(intermediate_reg_1[1417])); 
xor_module xor_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2833]),.i2(intermediate_reg_0[2832]),.o(intermediate_reg_1[1416])); 
mux_module mux_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2831]),.i2(intermediate_reg_0[2830]),.o(intermediate_reg_1[1415]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2829]),.i2(intermediate_reg_0[2828]),.o(intermediate_reg_1[1414])); 
xor_module xor_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2827]),.i2(intermediate_reg_0[2826]),.o(intermediate_reg_1[1413])); 
xor_module xor_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2825]),.i2(intermediate_reg_0[2824]),.o(intermediate_reg_1[1412])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2823]),.i2(intermediate_reg_0[2822]),.o(intermediate_reg_1[1411]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2821]),.i2(intermediate_reg_0[2820]),.o(intermediate_reg_1[1410]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2819]),.i2(intermediate_reg_0[2818]),.o(intermediate_reg_1[1409])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2817]),.i2(intermediate_reg_0[2816]),.o(intermediate_reg_1[1408])); 
xor_module xor_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2815]),.i2(intermediate_reg_0[2814]),.o(intermediate_reg_1[1407])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2813]),.i2(intermediate_reg_0[2812]),.o(intermediate_reg_1[1406])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2811]),.i2(intermediate_reg_0[2810]),.o(intermediate_reg_1[1405]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2809]),.i2(intermediate_reg_0[2808]),.o(intermediate_reg_1[1404])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2807]),.i2(intermediate_reg_0[2806]),.o(intermediate_reg_1[1403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2805]),.i2(intermediate_reg_0[2804]),.o(intermediate_reg_1[1402]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2803]),.i2(intermediate_reg_0[2802]),.o(intermediate_reg_1[1401]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2801]),.i2(intermediate_reg_0[2800]),.o(intermediate_reg_1[1400])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2799]),.i2(intermediate_reg_0[2798]),.o(intermediate_reg_1[1399]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2797]),.i2(intermediate_reg_0[2796]),.o(intermediate_reg_1[1398]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2795]),.i2(intermediate_reg_0[2794]),.o(intermediate_reg_1[1397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2793]),.i2(intermediate_reg_0[2792]),.o(intermediate_reg_1[1396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2791]),.i2(intermediate_reg_0[2790]),.o(intermediate_reg_1[1395])); 
xor_module xor_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2789]),.i2(intermediate_reg_0[2788]),.o(intermediate_reg_1[1394])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2787]),.i2(intermediate_reg_0[2786]),.o(intermediate_reg_1[1393])); 
mux_module mux_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2785]),.i2(intermediate_reg_0[2784]),.o(intermediate_reg_1[1392]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2783]),.i2(intermediate_reg_0[2782]),.o(intermediate_reg_1[1391])); 
mux_module mux_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2781]),.i2(intermediate_reg_0[2780]),.o(intermediate_reg_1[1390]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2779]),.i2(intermediate_reg_0[2778]),.o(intermediate_reg_1[1389]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2777]),.i2(intermediate_reg_0[2776]),.o(intermediate_reg_1[1388])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2775]),.i2(intermediate_reg_0[2774]),.o(intermediate_reg_1[1387]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2773]),.i2(intermediate_reg_0[2772]),.o(intermediate_reg_1[1386])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2771]),.i2(intermediate_reg_0[2770]),.o(intermediate_reg_1[1385]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2769]),.i2(intermediate_reg_0[2768]),.o(intermediate_reg_1[1384])); 
xor_module xor_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2767]),.i2(intermediate_reg_0[2766]),.o(intermediate_reg_1[1383])); 
xor_module xor_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2765]),.i2(intermediate_reg_0[2764]),.o(intermediate_reg_1[1382])); 
xor_module xor_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2763]),.i2(intermediate_reg_0[2762]),.o(intermediate_reg_1[1381])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2761]),.i2(intermediate_reg_0[2760]),.o(intermediate_reg_1[1380]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2759]),.i2(intermediate_reg_0[2758]),.o(intermediate_reg_1[1379]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2757]),.i2(intermediate_reg_0[2756]),.o(intermediate_reg_1[1378])); 
xor_module xor_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2755]),.i2(intermediate_reg_0[2754]),.o(intermediate_reg_1[1377])); 
mux_module mux_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2753]),.i2(intermediate_reg_0[2752]),.o(intermediate_reg_1[1376]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2751]),.i2(intermediate_reg_0[2750]),.o(intermediate_reg_1[1375])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2749]),.i2(intermediate_reg_0[2748]),.o(intermediate_reg_1[1374]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2747]),.i2(intermediate_reg_0[2746]),.o(intermediate_reg_1[1373])); 
xor_module xor_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2745]),.i2(intermediate_reg_0[2744]),.o(intermediate_reg_1[1372])); 
mux_module mux_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2743]),.i2(intermediate_reg_0[2742]),.o(intermediate_reg_1[1371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2741]),.i2(intermediate_reg_0[2740]),.o(intermediate_reg_1[1370]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2739]),.i2(intermediate_reg_0[2738]),.o(intermediate_reg_1[1369]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2737]),.i2(intermediate_reg_0[2736]),.o(intermediate_reg_1[1368]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2735]),.i2(intermediate_reg_0[2734]),.o(intermediate_reg_1[1367]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2733]),.i2(intermediate_reg_0[2732]),.o(intermediate_reg_1[1366])); 
xor_module xor_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2731]),.i2(intermediate_reg_0[2730]),.o(intermediate_reg_1[1365])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2729]),.i2(intermediate_reg_0[2728]),.o(intermediate_reg_1[1364]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2727]),.i2(intermediate_reg_0[2726]),.o(intermediate_reg_1[1363])); 
mux_module mux_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2725]),.i2(intermediate_reg_0[2724]),.o(intermediate_reg_1[1362]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2723]),.i2(intermediate_reg_0[2722]),.o(intermediate_reg_1[1361])); 
xor_module xor_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2721]),.i2(intermediate_reg_0[2720]),.o(intermediate_reg_1[1360])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2719]),.i2(intermediate_reg_0[2718]),.o(intermediate_reg_1[1359]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2717]),.i2(intermediate_reg_0[2716]),.o(intermediate_reg_1[1358])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2715]),.i2(intermediate_reg_0[2714]),.o(intermediate_reg_1[1357]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2713]),.i2(intermediate_reg_0[2712]),.o(intermediate_reg_1[1356])); 
xor_module xor_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2711]),.i2(intermediate_reg_0[2710]),.o(intermediate_reg_1[1355])); 
mux_module mux_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2709]),.i2(intermediate_reg_0[2708]),.o(intermediate_reg_1[1354]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2707]),.i2(intermediate_reg_0[2706]),.o(intermediate_reg_1[1353])); 
mux_module mux_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2705]),.i2(intermediate_reg_0[2704]),.o(intermediate_reg_1[1352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2703]),.i2(intermediate_reg_0[2702]),.o(intermediate_reg_1[1351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2701]),.i2(intermediate_reg_0[2700]),.o(intermediate_reg_1[1350]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2699]),.i2(intermediate_reg_0[2698]),.o(intermediate_reg_1[1349])); 
xor_module xor_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2697]),.i2(intermediate_reg_0[2696]),.o(intermediate_reg_1[1348])); 
mux_module mux_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2695]),.i2(intermediate_reg_0[2694]),.o(intermediate_reg_1[1347]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2693]),.i2(intermediate_reg_0[2692]),.o(intermediate_reg_1[1346]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2691]),.i2(intermediate_reg_0[2690]),.o(intermediate_reg_1[1345]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2689]),.i2(intermediate_reg_0[2688]),.o(intermediate_reg_1[1344]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343])); 
xor_module xor_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342])); 
mux_module mux_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334])); 
xor_module xor_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333])); 
xor_module xor_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322])); 
mux_module mux_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318])); 
xor_module xor_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315])); 
mux_module mux_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311])); 
xor_module xor_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310])); 
mux_module mux_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303])); 
mux_module mux_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301])); 
xor_module xor_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300])); 
mux_module mux_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298])); 
xor_module xor_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297])); 
mux_module mux_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294])); 
mux_module mux_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292])); 
xor_module xor_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291])); 
mux_module mux_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289])); 
xor_module xor_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288])); 
mux_module mux_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286])); 
xor_module xor_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284])); 
mux_module mux_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282])); 
mux_module mux_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276])); 
mux_module mux_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274])); 
xor_module xor_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264])); 
mux_module mux_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262])); 
xor_module xor_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261])); 
mux_module mux_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253])); 
xor_module xor_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252])); 
xor_module xor_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248])); 
xor_module xor_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247])); 
mux_module mux_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245])); 
mux_module mux_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241])); 
xor_module xor_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239])); 
xor_module xor_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238])); 
xor_module xor_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237])); 
xor_module xor_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236])); 
xor_module xor_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235])); 
xor_module xor_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234])); 
mux_module mux_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231])); 
mux_module mux_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228])); 
mux_module mux_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
mux_module mux_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222])); 
xor_module xor_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
mux_module mux_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219])); 
mux_module mux_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217])); 
xor_module xor_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216])); 
xor_module xor_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215])); 
xor_module xor_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209])); 
mux_module mux_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207])); 
mux_module mux_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205])); 
xor_module xor_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198])); 
xor_module xor_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197])); 
xor_module xor_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196])); 
xor_module xor_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195])); 
mux_module mux_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193])); 
mux_module mux_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191])); 
xor_module xor_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187])); 
mux_module mux_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184])); 
xor_module xor_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183])); 
xor_module xor_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182])); 
xor_module xor_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181])); 
mux_module mux_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179])); 
xor_module xor_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178])); 
xor_module xor_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177])); 
xor_module xor_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176])); 
mux_module mux_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174])); 
mux_module mux_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172])); 
mux_module mux_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161])); 
mux_module mux_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
mux_module mux_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155])); 
xor_module xor_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154])); 
xor_module xor_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153])); 
mux_module mux_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151])); 
mux_module mux_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149])); 
mux_module mux_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146])); 
mux_module mux_module_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142])); 
mux_module mux_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140])); 
mux_module mux_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138])); 
xor_module xor_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137])); 
xor_module xor_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136])); 
xor_module xor_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135])); 
xor_module xor_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134])); 
mux_module mux_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132])); 
mux_module mux_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
xor_module xor_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129])); 
mux_module mux_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127])); 
mux_module mux_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
xor_module xor_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
xor_module xor_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123])); 
mux_module mux_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120])); 
xor_module xor_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
mux_module mux_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114])); 
xor_module xor_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113])); 
xor_module xor_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112])); 
xor_module xor_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111])); 
xor_module xor_module_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110])); 
xor_module xor_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109])); 
xor_module xor_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
mux_module mux_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
mux_module mux_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102])); 
xor_module xor_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
mux_module mux_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097])); 
xor_module xor_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096])); 
xor_module xor_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095])); 
xor_module xor_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094])); 
mux_module mux_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
mux_module mux_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090])); 
xor_module xor_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
xor_module xor_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086])); 
xor_module xor_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085])); 
mux_module mux_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082])); 
mux_module mux_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080])); 
xor_module xor_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079])); 
mux_module mux_module_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076])); 
mux_module mux_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074])); 
xor_module xor_module_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
mux_module mux_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071])); 
mux_module mux_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069])); 
xor_module xor_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068])); 
xor_module xor_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
xor_module xor_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066])); 
xor_module xor_module_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065])); 
xor_module xor_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064])); 
mux_module mux_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062])); 
mux_module mux_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056])); 
xor_module xor_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053])); 
xor_module xor_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
xor_module xor_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051])); 
xor_module xor_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050])); 
xor_module xor_module_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049])); 
mux_module mux_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
mux_module mux_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038])); 
mux_module mux_module_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036])); 
xor_module xor_module_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035])); 
xor_module xor_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034])); 
xor_module xor_module_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033])); 
mux_module mux_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030])); 
mux_module mux_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
mux_module mux_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
xor_module xor_module_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022])); 
xor_module xor_module_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021])); 
xor_module xor_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
mux_module mux_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018])); 
mux_module mux_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016])); 
xor_module xor_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
xor_module xor_module_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
mux_module mux_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
xor_module xor_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
mux_module mux_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
mux_module mux_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
xor_module xor_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999])); 
xor_module xor_module_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
mux_module mux_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
xor_module xor_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
xor_module xor_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
xor_module xor_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
mux_module mux_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
mux_module mux_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
mux_module mux_module_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
mux_module mux_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
xor_module xor_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
mux_module mux_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
xor_module xor_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
mux_module mux_module_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
xor_module xor_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962])); 
mux_module mux_module_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
mux_module mux_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
mux_module mux_module_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
xor_module xor_module_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
mux_module mux_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948])); 
mux_module mux_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
xor_module xor_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
xor_module xor_module_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
xor_module xor_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
xor_module xor_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
xor_module xor_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
mux_module mux_module_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
mux_module mux_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
mux_module mux_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
mux_module mux_module_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
xor_module xor_module_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
xor_module xor_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
mux_module mux_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
mux_module mux_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
xor_module xor_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
mux_module mux_module_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
xor_module xor_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
xor_module xor_module_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
xor_module xor_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
xor_module xor_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
xor_module xor_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
xor_module xor_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
mux_module mux_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
mux_module mux_module_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906])); 
xor_module xor_module_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
xor_module xor_module_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
xor_module xor_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
mux_module mux_module_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
xor_module xor_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
mux_module mux_module_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
mux_module mux_module_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
xor_module xor_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
mux_module mux_module_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
mux_module mux_module_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
mux_module mux_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
mux_module mux_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879])); 
mux_module mux_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
mux_module mux_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
xor_module xor_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
mux_module mux_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
mux_module mux_module_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
xor_module xor_module_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
mux_module mux_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
mux_module mux_module_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862])); 
mux_module mux_module_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
mux_module mux_module_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
mux_module mux_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
xor_module xor_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
xor_module xor_module_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
mux_module mux_module_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
mux_module mux_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
xor_module xor_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
xor_module xor_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
xor_module xor_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
mux_module mux_module_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
xor_module xor_module_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
mux_module mux_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829])); 
mux_module mux_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
xor_module xor_module_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
xor_module xor_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823])); 
xor_module xor_module_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
mux_module mux_module_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
mux_module mux_module_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
xor_module xor_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
mux_module mux_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
mux_module mux_module_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
xor_module xor_module_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
xor_module xor_module_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
mux_module mux_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
xor_module xor_module_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
xor_module xor_module_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
xor_module xor_module_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
mux_module mux_module_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
xor_module xor_module_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
mux_module mux_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
xor_module xor_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
mux_module mux_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
mux_module mux_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
xor_module xor_module_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
xor_module xor_module_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
xor_module xor_module_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
mux_module mux_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
mux_module mux_module_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
xor_module xor_module_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
xor_module xor_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
xor_module xor_module_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
mux_module mux_module_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
xor_module xor_module_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
xor_module xor_module_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
mux_module mux_module_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
xor_module xor_module_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
mux_module mux_module_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
xor_module xor_module_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
xor_module xor_module_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
xor_module xor_module_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
xor_module xor_module_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
xor_module xor_module_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
mux_module mux_module_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
xor_module xor_module_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
xor_module xor_module_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
mux_module mux_module_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
mux_module mux_module_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
mux_module mux_module_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
xor_module xor_module_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
mux_module mux_module_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
mux_module mux_module_inst_1_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
mux_module mux_module_inst_1_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
mux_module mux_module_inst_1_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
xor_module xor_module_inst_1_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
mux_module mux_module_inst_1_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
xor_module xor_module_inst_1_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
xor_module xor_module_inst_1_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
mux_module mux_module_inst_1_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
mux_module mux_module_inst_1_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
xor_module xor_module_inst_1_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
mux_module mux_module_inst_1_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
mux_module mux_module_inst_1_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
mux_module mux_module_inst_1_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
mux_module mux_module_inst_1_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
mux_module mux_module_inst_1_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
mux_module mux_module_inst_1_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
mux_module mux_module_inst_1_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
xor_module xor_module_inst_1_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
xor_module xor_module_inst_1_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
xor_module xor_module_inst_1_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
mux_module mux_module_inst_1_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
xor_module xor_module_inst_1_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
mux_module mux_module_inst_1_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
mux_module mux_module_inst_1_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
xor_module xor_module_inst_1_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
mux_module mux_module_inst_1_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
mux_module mux_module_inst_1_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
mux_module mux_module_inst_1_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
xor_module xor_module_inst_1_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
mux_module mux_module_inst_1_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
mux_module mux_module_inst_1_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
mux_module mux_module_inst_1_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
xor_module xor_module_inst_1_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
mux_module mux_module_inst_1_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
mux_module mux_module_inst_1_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
mux_module mux_module_inst_1_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
xor_module xor_module_inst_1_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
xor_module xor_module_inst_1_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
mux_module mux_module_inst_1_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
mux_module mux_module_inst_1_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
xor_module xor_module_inst_1_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
xor_module xor_module_inst_1_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
xor_module xor_module_inst_1_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
mux_module mux_module_inst_1_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
xor_module xor_module_inst_1_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
mux_module mux_module_inst_1_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
xor_module xor_module_inst_1_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
xor_module xor_module_inst_1_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
mux_module mux_module_inst_1_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
xor_module xor_module_inst_1_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
xor_module xor_module_inst_1_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
mux_module mux_module_inst_1_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
mux_module mux_module_inst_1_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
xor_module xor_module_inst_1_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
xor_module xor_module_inst_1_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
xor_module xor_module_inst_1_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
xor_module xor_module_inst_1_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
mux_module mux_module_inst_1_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
mux_module mux_module_inst_1_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
xor_module xor_module_inst_1_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
mux_module mux_module_inst_1_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
xor_module xor_module_inst_1_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
xor_module xor_module_inst_1_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
mux_module mux_module_inst_1_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
xor_module xor_module_inst_1_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
mux_module mux_module_inst_1_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
xor_module xor_module_inst_1_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
mux_module mux_module_inst_1_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
mux_module mux_module_inst_1_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
xor_module xor_module_inst_1_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
mux_module mux_module_inst_1_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
xor_module xor_module_inst_1_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
xor_module xor_module_inst_1_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
xor_module xor_module_inst_1_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
mux_module mux_module_inst_1_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
mux_module mux_module_inst_1_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
mux_module mux_module_inst_1_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
xor_module xor_module_inst_1_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
mux_module mux_module_inst_1_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
mux_module mux_module_inst_1_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
mux_module mux_module_inst_1_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
mux_module mux_module_inst_1_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
mux_module mux_module_inst_1_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
xor_module xor_module_inst_1_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
xor_module xor_module_inst_1_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
xor_module xor_module_inst_1_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
xor_module xor_module_inst_1_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
mux_module mux_module_inst_1_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
xor_module xor_module_inst_1_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
mux_module mux_module_inst_1_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
xor_module xor_module_inst_1_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
mux_module mux_module_inst_1_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
mux_module mux_module_inst_1_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
xor_module xor_module_inst_1_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
mux_module mux_module_inst_1_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
xor_module xor_module_inst_1_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
xor_module xor_module_inst_1_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
mux_module mux_module_inst_1_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
mux_module mux_module_inst_1_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
mux_module mux_module_inst_1_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
xor_module xor_module_inst_1_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
mux_module mux_module_inst_1_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
xor_module xor_module_inst_1_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
mux_module mux_module_inst_1_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
xor_module xor_module_inst_1_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
mux_module mux_module_inst_1_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
xor_module xor_module_inst_1_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
mux_module mux_module_inst_1_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
mux_module mux_module_inst_1_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
xor_module xor_module_inst_1_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
xor_module xor_module_inst_1_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
mux_module mux_module_inst_1_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
xor_module xor_module_inst_1_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
xor_module xor_module_inst_1_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
mux_module mux_module_inst_1_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
mux_module mux_module_inst_1_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
xor_module xor_module_inst_1_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
mux_module mux_module_inst_1_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
xor_module xor_module_inst_1_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
mux_module mux_module_inst_1_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
mux_module mux_module_inst_1_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
xor_module xor_module_inst_1_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
xor_module xor_module_inst_1_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
mux_module mux_module_inst_1_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
xor_module xor_module_inst_1_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
mux_module mux_module_inst_1_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
mux_module mux_module_inst_1_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
xor_module xor_module_inst_1_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
mux_module mux_module_inst_1_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
mux_module mux_module_inst_1_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
mux_module mux_module_inst_1_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
xor_module xor_module_inst_1_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
xor_module xor_module_inst_1_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
xor_module xor_module_inst_1_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
mux_module mux_module_inst_1_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
xor_module xor_module_inst_1_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
xor_module xor_module_inst_1_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
mux_module mux_module_inst_1_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
mux_module mux_module_inst_1_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
mux_module mux_module_inst_1_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
xor_module xor_module_inst_1_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
mux_module mux_module_inst_1_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
mux_module mux_module_inst_1_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
mux_module mux_module_inst_1_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
mux_module mux_module_inst_1_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
mux_module mux_module_inst_1_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
mux_module mux_module_inst_1_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
mux_module mux_module_inst_1_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
xor_module xor_module_inst_1_1650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
mux_module mux_module_inst_1_1651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
mux_module mux_module_inst_1_1655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
xor_module xor_module_inst_1_1658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
xor_module xor_module_inst_1_1659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
xor_module xor_module_inst_1_1660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
mux_module mux_module_inst_1_1661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
mux_module mux_module_inst_1_1663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
mux_module mux_module_inst_1_1665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_1668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
xor_module xor_module_inst_1_1669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
mux_module mux_module_inst_1_1670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
mux_module mux_module_inst_1_1674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
mux_module mux_module_inst_1_1676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_1679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
xor_module xor_module_inst_1_1681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
mux_module mux_module_inst_1_1682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
xor_module xor_module_inst_1_1684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
mux_module mux_module_inst_1_1685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
mux_module mux_module_inst_1_1689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
xor_module xor_module_inst_1_1691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
mux_module mux_module_inst_1_1692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
xor_module xor_module_inst_1_1695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_1696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
mux_module mux_module_inst_1_1698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
mux_module mux_module_inst_1_1703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
mux_module mux_module_inst_1_1711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
xor_module xor_module_inst_1_1713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
mux_module mux_module_inst_1_1714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
xor_module xor_module_inst_1_1716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
mux_module mux_module_inst_1_1717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
mux_module mux_module_inst_1_1719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
mux_module mux_module_inst_1_1722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
xor_module xor_module_inst_1_1725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
mux_module mux_module_inst_1_1726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
xor_module xor_module_inst_1_1729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
mux_module mux_module_inst_1_1730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
mux_module mux_module_inst_1_1735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
xor_module xor_module_inst_1_1737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
xor_module xor_module_inst_1_1738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
mux_module mux_module_inst_1_1739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_1741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
xor_module xor_module_inst_1_1746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
mux_module mux_module_inst_1_1747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
mux_module mux_module_inst_1_1749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
xor_module xor_module_inst_1_1752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
mux_module mux_module_inst_1_1753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
xor_module xor_module_inst_1_1757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
mux_module mux_module_inst_1_1758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
xor_module xor_module_inst_1_1762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
mux_module mux_module_inst_1_1763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
xor_module xor_module_inst_1_1765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
xor_module xor_module_inst_1_1766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
mux_module mux_module_inst_1_1767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
xor_module xor_module_inst_1_1770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
mux_module mux_module_inst_1_1771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
mux_module mux_module_inst_1_1773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
mux_module mux_module_inst_1_1775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
mux_module mux_module_inst_1_1777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
xor_module xor_module_inst_1_1779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
mux_module mux_module_inst_1_1780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
mux_module mux_module_inst_1_1782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
xor_module xor_module_inst_1_1787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
mux_module mux_module_inst_1_1788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
xor_module xor_module_inst_1_1791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
mux_module mux_module_inst_1_1792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
mux_module mux_module_inst_1_1795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
mux_module mux_module_inst_1_1797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
mux_module mux_module_inst_1_1799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
xor_module xor_module_inst_1_1802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
xor_module xor_module_inst_1_1803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
mux_module mux_module_inst_1_1804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
xor_module xor_module_inst_1_1806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
mux_module mux_module_inst_1_1807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
mux_module mux_module_inst_1_1813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
mux_module mux_module_inst_1_1816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
xor_module xor_module_inst_1_1822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
xor_module xor_module_inst_1_1823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
mux_module mux_module_inst_1_1824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
mux_module mux_module_inst_1_1827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
mux_module mux_module_inst_1_1829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
xor_module xor_module_inst_1_1831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
xor_module xor_module_inst_1_1832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
mux_module mux_module_inst_1_1833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
mux_module mux_module_inst_1_1836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
xor_module xor_module_inst_1_1839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
xor_module xor_module_inst_1_1840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
xor_module xor_module_inst_1_1841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_1842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
mux_module mux_module_inst_1_1843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
xor_module xor_module_inst_1_1850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
xor_module xor_module_inst_1_1851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
xor_module xor_module_inst_1_1852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
mux_module mux_module_inst_1_1853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
xor_module xor_module_inst_1_1857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
mux_module mux_module_inst_1_1858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
mux_module mux_module_inst_1_1861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
xor_module xor_module_inst_1_1863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
xor_module xor_module_inst_1_1864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
xor_module xor_module_inst_1_1865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
mux_module mux_module_inst_1_1866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
mux_module mux_module_inst_1_1870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_1873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_1874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
xor_module xor_module_inst_1_1878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
mux_module mux_module_inst_1_1879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
mux_module mux_module_inst_1_1881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
mux_module mux_module_inst_1_1884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
xor_module xor_module_inst_1_1886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
xor_module xor_module_inst_1_1887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
xor_module xor_module_inst_1_1888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
xor_module xor_module_inst_1_1889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
mux_module mux_module_inst_1_1890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
mux_module mux_module_inst_1_1892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
mux_module mux_module_inst_1_1894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
xor_module xor_module_inst_1_1896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
xor_module xor_module_inst_1_1897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
xor_module xor_module_inst_1_1898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
mux_module mux_module_inst_1_1899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
xor_module xor_module_inst_1_1902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
xor_module xor_module_inst_1_1903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
xor_module xor_module_inst_1_1904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
mux_module mux_module_inst_1_1905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
xor_module xor_module_inst_1_1908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
mux_module mux_module_inst_1_1909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
mux_module mux_module_inst_1_1917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
mux_module mux_module_inst_1_1923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
mux_module mux_module_inst_1_1925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
xor_module xor_module_inst_1_1929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
mux_module mux_module_inst_1_1930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
mux_module mux_module_inst_1_1933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
xor_module xor_module_inst_1_1936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
xor_module xor_module_inst_1_1937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
mux_module mux_module_inst_1_1938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
mux_module mux_module_inst_1_1944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
xor_module xor_module_inst_1_1948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
mux_module mux_module_inst_1_1949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
mux_module mux_module_inst_1_1951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
xor_module xor_module_inst_1_1953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_1954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_1955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
xor_module xor_module_inst_1_1956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_1957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
xor_module xor_module_inst_1_1958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
xor_module xor_module_inst_1_1959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
mux_module mux_module_inst_1_1960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
xor_module xor_module_inst_1_1962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
mux_module mux_module_inst_1_1963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
mux_module mux_module_inst_1_1965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
mux_module mux_module_inst_1_1967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
xor_module xor_module_inst_1_1972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
xor_module xor_module_inst_1_1973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
mux_module mux_module_inst_1_1974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
mux_module mux_module_inst_1_1980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
xor_module xor_module_inst_1_1985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
xor_module xor_module_inst_1_1986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
xor_module xor_module_inst_1_1987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
mux_module mux_module_inst_1_1988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
mux_module mux_module_inst_1_1990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
xor_module xor_module_inst_1_1992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
xor_module xor_module_inst_1_1993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
xor_module xor_module_inst_1_1994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
xor_module xor_module_inst_1_1995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_1996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_1997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
mux_module mux_module_inst_1_1998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_2000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
xor_module xor_module_inst_1_2001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
xor_module xor_module_inst_1_2002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
xor_module xor_module_inst_1_2003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
mux_module mux_module_inst_1_2004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
xor_module xor_module_inst_1_2006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
mux_module mux_module_inst_1_2007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_2009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
mux_module mux_module_inst_1_2012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
xor_module xor_module_inst_1_2014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
mux_module mux_module_inst_1_2015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
mux_module mux_module_inst_1_2021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
mux_module mux_module_inst_1_2027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
xor_module xor_module_inst_1_2029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
xor_module xor_module_inst_1_2030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
xor_module xor_module_inst_1_2031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
mux_module mux_module_inst_1_2032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
xor_module xor_module_inst_1_2036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
xor_module xor_module_inst_1_2037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
mux_module mux_module_inst_1_2038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_2041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
mux_module mux_module_inst_1_2042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
xor_module xor_module_inst_1_2045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
mux_module mux_module_inst_1_2046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
xor_module xor_module_inst_1_2048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_2049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
mux_module mux_module_inst_1_2050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
mux_module mux_module_inst_1_2054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_2057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_2059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_2060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
xor_module xor_module_inst_1_2061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
xor_module xor_module_inst_1_2062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
xor_module xor_module_inst_1_2063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
mux_module mux_module_inst_1_2064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_2068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
xor_module xor_module_inst_1_2069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
xor_module xor_module_inst_1_2070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
xor_module xor_module_inst_1_2071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
reg [1035:0]intermediate_reg_2; 
 
xor_module xor_module_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2071]),.i2(intermediate_reg_1[2070]),.o(intermediate_reg_2[1035])); 
xor_module xor_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2069]),.i2(intermediate_reg_1[2068]),.o(intermediate_reg_2[1034])); 
xor_module xor_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2067]),.i2(intermediate_reg_1[2066]),.o(intermediate_reg_2[1033])); 
xor_module xor_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2065]),.i2(intermediate_reg_1[2064]),.o(intermediate_reg_2[1032])); 
mux_module mux_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2063]),.i2(intermediate_reg_1[2062]),.o(intermediate_reg_2[1031]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2061]),.i2(intermediate_reg_1[2060]),.o(intermediate_reg_2[1030])); 
mux_module mux_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2059]),.i2(intermediate_reg_1[2058]),.o(intermediate_reg_2[1029]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2057]),.i2(intermediate_reg_1[2056]),.o(intermediate_reg_2[1028])); 
xor_module xor_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2055]),.i2(intermediate_reg_1[2054]),.o(intermediate_reg_2[1027])); 
mux_module mux_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2053]),.i2(intermediate_reg_1[2052]),.o(intermediate_reg_2[1026]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2051]),.i2(intermediate_reg_1[2050]),.o(intermediate_reg_2[1025]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2049]),.i2(intermediate_reg_1[2048]),.o(intermediate_reg_2[1024]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2047]),.i2(intermediate_reg_1[2046]),.o(intermediate_reg_2[1023])); 
mux_module mux_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2045]),.i2(intermediate_reg_1[2044]),.o(intermediate_reg_2[1022]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2043]),.i2(intermediate_reg_1[2042]),.o(intermediate_reg_2[1021])); 
mux_module mux_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2041]),.i2(intermediate_reg_1[2040]),.o(intermediate_reg_2[1020]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2039]),.i2(intermediate_reg_1[2038]),.o(intermediate_reg_2[1019])); 
mux_module mux_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2037]),.i2(intermediate_reg_1[2036]),.o(intermediate_reg_2[1018]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2035]),.i2(intermediate_reg_1[2034]),.o(intermediate_reg_2[1017]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2033]),.i2(intermediate_reg_1[2032]),.o(intermediate_reg_2[1016])); 
xor_module xor_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2031]),.i2(intermediate_reg_1[2030]),.o(intermediate_reg_2[1015])); 
mux_module mux_module_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2029]),.i2(intermediate_reg_1[2028]),.o(intermediate_reg_2[1014]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2027]),.i2(intermediate_reg_1[2026]),.o(intermediate_reg_2[1013]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2025]),.i2(intermediate_reg_1[2024]),.o(intermediate_reg_2[1012]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2023]),.i2(intermediate_reg_1[2022]),.o(intermediate_reg_2[1011]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2021]),.i2(intermediate_reg_1[2020]),.o(intermediate_reg_2[1010]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2019]),.i2(intermediate_reg_1[2018]),.o(intermediate_reg_2[1009])); 
mux_module mux_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2017]),.i2(intermediate_reg_1[2016]),.o(intermediate_reg_2[1008]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2015]),.i2(intermediate_reg_1[2014]),.o(intermediate_reg_2[1007]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2013]),.i2(intermediate_reg_1[2012]),.o(intermediate_reg_2[1006]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2011]),.i2(intermediate_reg_1[2010]),.o(intermediate_reg_2[1005])); 
xor_module xor_module_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2009]),.i2(intermediate_reg_1[2008]),.o(intermediate_reg_2[1004])); 
mux_module mux_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2007]),.i2(intermediate_reg_1[2006]),.o(intermediate_reg_2[1003]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2005]),.i2(intermediate_reg_1[2004]),.o(intermediate_reg_2[1002])); 
mux_module mux_module_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2003]),.i2(intermediate_reg_1[2002]),.o(intermediate_reg_2[1001]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[2001]),.i2(intermediate_reg_1[2000]),.o(intermediate_reg_2[1000]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1999]),.i2(intermediate_reg_1[1998]),.o(intermediate_reg_2[999]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1997]),.i2(intermediate_reg_1[1996]),.o(intermediate_reg_2[998]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1995]),.i2(intermediate_reg_1[1994]),.o(intermediate_reg_2[997]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1993]),.i2(intermediate_reg_1[1992]),.o(intermediate_reg_2[996]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1991]),.i2(intermediate_reg_1[1990]),.o(intermediate_reg_2[995]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1989]),.i2(intermediate_reg_1[1988]),.o(intermediate_reg_2[994])); 
mux_module mux_module_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1987]),.i2(intermediate_reg_1[1986]),.o(intermediate_reg_2[993]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1985]),.i2(intermediate_reg_1[1984]),.o(intermediate_reg_2[992]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1983]),.i2(intermediate_reg_1[1982]),.o(intermediate_reg_2[991]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1981]),.i2(intermediate_reg_1[1980]),.o(intermediate_reg_2[990]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1979]),.i2(intermediate_reg_1[1978]),.o(intermediate_reg_2[989])); 
mux_module mux_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1977]),.i2(intermediate_reg_1[1976]),.o(intermediate_reg_2[988]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1975]),.i2(intermediate_reg_1[1974]),.o(intermediate_reg_2[987]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1973]),.i2(intermediate_reg_1[1972]),.o(intermediate_reg_2[986])); 
xor_module xor_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1971]),.i2(intermediate_reg_1[1970]),.o(intermediate_reg_2[985])); 
mux_module mux_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1969]),.i2(intermediate_reg_1[1968]),.o(intermediate_reg_2[984]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1967]),.i2(intermediate_reg_1[1966]),.o(intermediate_reg_2[983])); 
xor_module xor_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1965]),.i2(intermediate_reg_1[1964]),.o(intermediate_reg_2[982])); 
xor_module xor_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1963]),.i2(intermediate_reg_1[1962]),.o(intermediate_reg_2[981])); 
xor_module xor_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1961]),.i2(intermediate_reg_1[1960]),.o(intermediate_reg_2[980])); 
xor_module xor_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1959]),.i2(intermediate_reg_1[1958]),.o(intermediate_reg_2[979])); 
xor_module xor_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1957]),.i2(intermediate_reg_1[1956]),.o(intermediate_reg_2[978])); 
mux_module mux_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1955]),.i2(intermediate_reg_1[1954]),.o(intermediate_reg_2[977]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1953]),.i2(intermediate_reg_1[1952]),.o(intermediate_reg_2[976])); 
mux_module mux_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1951]),.i2(intermediate_reg_1[1950]),.o(intermediate_reg_2[975]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1949]),.i2(intermediate_reg_1[1948]),.o(intermediate_reg_2[974])); 
xor_module xor_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1947]),.i2(intermediate_reg_1[1946]),.o(intermediate_reg_2[973])); 
mux_module mux_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1945]),.i2(intermediate_reg_1[1944]),.o(intermediate_reg_2[972]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1943]),.i2(intermediate_reg_1[1942]),.o(intermediate_reg_2[971])); 
mux_module mux_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1941]),.i2(intermediate_reg_1[1940]),.o(intermediate_reg_2[970]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1939]),.i2(intermediate_reg_1[1938]),.o(intermediate_reg_2[969])); 
mux_module mux_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1937]),.i2(intermediate_reg_1[1936]),.o(intermediate_reg_2[968]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1935]),.i2(intermediate_reg_1[1934]),.o(intermediate_reg_2[967]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1933]),.i2(intermediate_reg_1[1932]),.o(intermediate_reg_2[966])); 
mux_module mux_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1931]),.i2(intermediate_reg_1[1930]),.o(intermediate_reg_2[965]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1929]),.i2(intermediate_reg_1[1928]),.o(intermediate_reg_2[964]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1927]),.i2(intermediate_reg_1[1926]),.o(intermediate_reg_2[963]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1925]),.i2(intermediate_reg_1[1924]),.o(intermediate_reg_2[962])); 
xor_module xor_module_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1923]),.i2(intermediate_reg_1[1922]),.o(intermediate_reg_2[961])); 
xor_module xor_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1921]),.i2(intermediate_reg_1[1920]),.o(intermediate_reg_2[960])); 
xor_module xor_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1919]),.i2(intermediate_reg_1[1918]),.o(intermediate_reg_2[959])); 
mux_module mux_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1917]),.i2(intermediate_reg_1[1916]),.o(intermediate_reg_2[958]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1915]),.i2(intermediate_reg_1[1914]),.o(intermediate_reg_2[957]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1913]),.i2(intermediate_reg_1[1912]),.o(intermediate_reg_2[956])); 
mux_module mux_module_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1911]),.i2(intermediate_reg_1[1910]),.o(intermediate_reg_2[955]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1909]),.i2(intermediate_reg_1[1908]),.o(intermediate_reg_2[954])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1907]),.i2(intermediate_reg_1[1906]),.o(intermediate_reg_2[953]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1905]),.i2(intermediate_reg_1[1904]),.o(intermediate_reg_2[952]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1903]),.i2(intermediate_reg_1[1902]),.o(intermediate_reg_2[951]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1901]),.i2(intermediate_reg_1[1900]),.o(intermediate_reg_2[950]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1899]),.i2(intermediate_reg_1[1898]),.o(intermediate_reg_2[949])); 
xor_module xor_module_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1897]),.i2(intermediate_reg_1[1896]),.o(intermediate_reg_2[948])); 
mux_module mux_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1895]),.i2(intermediate_reg_1[1894]),.o(intermediate_reg_2[947]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1893]),.i2(intermediate_reg_1[1892]),.o(intermediate_reg_2[946])); 
xor_module xor_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1891]),.i2(intermediate_reg_1[1890]),.o(intermediate_reg_2[945])); 
mux_module mux_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1889]),.i2(intermediate_reg_1[1888]),.o(intermediate_reg_2[944]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1887]),.i2(intermediate_reg_1[1886]),.o(intermediate_reg_2[943]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1885]),.i2(intermediate_reg_1[1884]),.o(intermediate_reg_2[942]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1883]),.i2(intermediate_reg_1[1882]),.o(intermediate_reg_2[941])); 
mux_module mux_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1881]),.i2(intermediate_reg_1[1880]),.o(intermediate_reg_2[940]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1879]),.i2(intermediate_reg_1[1878]),.o(intermediate_reg_2[939])); 
xor_module xor_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1877]),.i2(intermediate_reg_1[1876]),.o(intermediate_reg_2[938])); 
xor_module xor_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1875]),.i2(intermediate_reg_1[1874]),.o(intermediate_reg_2[937])); 
xor_module xor_module_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1873]),.i2(intermediate_reg_1[1872]),.o(intermediate_reg_2[936])); 
xor_module xor_module_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1871]),.i2(intermediate_reg_1[1870]),.o(intermediate_reg_2[935])); 
mux_module mux_module_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1869]),.i2(intermediate_reg_1[1868]),.o(intermediate_reg_2[934]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1867]),.i2(intermediate_reg_1[1866]),.o(intermediate_reg_2[933])); 
mux_module mux_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1865]),.i2(intermediate_reg_1[1864]),.o(intermediate_reg_2[932]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1863]),.i2(intermediate_reg_1[1862]),.o(intermediate_reg_2[931])); 
xor_module xor_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1861]),.i2(intermediate_reg_1[1860]),.o(intermediate_reg_2[930])); 
mux_module mux_module_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1859]),.i2(intermediate_reg_1[1858]),.o(intermediate_reg_2[929]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1857]),.i2(intermediate_reg_1[1856]),.o(intermediate_reg_2[928])); 
mux_module mux_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1855]),.i2(intermediate_reg_1[1854]),.o(intermediate_reg_2[927]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1853]),.i2(intermediate_reg_1[1852]),.o(intermediate_reg_2[926])); 
xor_module xor_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1851]),.i2(intermediate_reg_1[1850]),.o(intermediate_reg_2[925])); 
xor_module xor_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1849]),.i2(intermediate_reg_1[1848]),.o(intermediate_reg_2[924])); 
mux_module mux_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1847]),.i2(intermediate_reg_1[1846]),.o(intermediate_reg_2[923]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1845]),.i2(intermediate_reg_1[1844]),.o(intermediate_reg_2[922]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1843]),.i2(intermediate_reg_1[1842]),.o(intermediate_reg_2[921])); 
xor_module xor_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1841]),.i2(intermediate_reg_1[1840]),.o(intermediate_reg_2[920])); 
mux_module mux_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1839]),.i2(intermediate_reg_1[1838]),.o(intermediate_reg_2[919]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1837]),.i2(intermediate_reg_1[1836]),.o(intermediate_reg_2[918])); 
mux_module mux_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1835]),.i2(intermediate_reg_1[1834]),.o(intermediate_reg_2[917]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1833]),.i2(intermediate_reg_1[1832]),.o(intermediate_reg_2[916]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1831]),.i2(intermediate_reg_1[1830]),.o(intermediate_reg_2[915])); 
xor_module xor_module_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1829]),.i2(intermediate_reg_1[1828]),.o(intermediate_reg_2[914])); 
mux_module mux_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1827]),.i2(intermediate_reg_1[1826]),.o(intermediate_reg_2[913]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1825]),.i2(intermediate_reg_1[1824]),.o(intermediate_reg_2[912])); 
mux_module mux_module_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1823]),.i2(intermediate_reg_1[1822]),.o(intermediate_reg_2[911]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1821]),.i2(intermediate_reg_1[1820]),.o(intermediate_reg_2[910])); 
xor_module xor_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1819]),.i2(intermediate_reg_1[1818]),.o(intermediate_reg_2[909])); 
mux_module mux_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1817]),.i2(intermediate_reg_1[1816]),.o(intermediate_reg_2[908]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1815]),.i2(intermediate_reg_1[1814]),.o(intermediate_reg_2[907])); 
xor_module xor_module_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1813]),.i2(intermediate_reg_1[1812]),.o(intermediate_reg_2[906])); 
xor_module xor_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1811]),.i2(intermediate_reg_1[1810]),.o(intermediate_reg_2[905])); 
mux_module mux_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1809]),.i2(intermediate_reg_1[1808]),.o(intermediate_reg_2[904]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1807]),.i2(intermediate_reg_1[1806]),.o(intermediate_reg_2[903]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1805]),.i2(intermediate_reg_1[1804]),.o(intermediate_reg_2[902]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1803]),.i2(intermediate_reg_1[1802]),.o(intermediate_reg_2[901]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1801]),.i2(intermediate_reg_1[1800]),.o(intermediate_reg_2[900]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1799]),.i2(intermediate_reg_1[1798]),.o(intermediate_reg_2[899]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1797]),.i2(intermediate_reg_1[1796]),.o(intermediate_reg_2[898])); 
mux_module mux_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1795]),.i2(intermediate_reg_1[1794]),.o(intermediate_reg_2[897]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1793]),.i2(intermediate_reg_1[1792]),.o(intermediate_reg_2[896])); 
xor_module xor_module_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1791]),.i2(intermediate_reg_1[1790]),.o(intermediate_reg_2[895])); 
mux_module mux_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1789]),.i2(intermediate_reg_1[1788]),.o(intermediate_reg_2[894]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1787]),.i2(intermediate_reg_1[1786]),.o(intermediate_reg_2[893])); 
xor_module xor_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1785]),.i2(intermediate_reg_1[1784]),.o(intermediate_reg_2[892])); 
mux_module mux_module_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1783]),.i2(intermediate_reg_1[1782]),.o(intermediate_reg_2[891]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1781]),.i2(intermediate_reg_1[1780]),.o(intermediate_reg_2[890]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1779]),.i2(intermediate_reg_1[1778]),.o(intermediate_reg_2[889]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1777]),.i2(intermediate_reg_1[1776]),.o(intermediate_reg_2[888])); 
xor_module xor_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1775]),.i2(intermediate_reg_1[1774]),.o(intermediate_reg_2[887])); 
xor_module xor_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1773]),.i2(intermediate_reg_1[1772]),.o(intermediate_reg_2[886])); 
mux_module mux_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1771]),.i2(intermediate_reg_1[1770]),.o(intermediate_reg_2[885]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1769]),.i2(intermediate_reg_1[1768]),.o(intermediate_reg_2[884]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1767]),.i2(intermediate_reg_1[1766]),.o(intermediate_reg_2[883])); 
mux_module mux_module_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1765]),.i2(intermediate_reg_1[1764]),.o(intermediate_reg_2[882]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1763]),.i2(intermediate_reg_1[1762]),.o(intermediate_reg_2[881])); 
mux_module mux_module_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1761]),.i2(intermediate_reg_1[1760]),.o(intermediate_reg_2[880]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1759]),.i2(intermediate_reg_1[1758]),.o(intermediate_reg_2[879]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1757]),.i2(intermediate_reg_1[1756]),.o(intermediate_reg_2[878]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1755]),.i2(intermediate_reg_1[1754]),.o(intermediate_reg_2[877]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1753]),.i2(intermediate_reg_1[1752]),.o(intermediate_reg_2[876]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1751]),.i2(intermediate_reg_1[1750]),.o(intermediate_reg_2[875])); 
xor_module xor_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1749]),.i2(intermediate_reg_1[1748]),.o(intermediate_reg_2[874])); 
xor_module xor_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1747]),.i2(intermediate_reg_1[1746]),.o(intermediate_reg_2[873])); 
mux_module mux_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1745]),.i2(intermediate_reg_1[1744]),.o(intermediate_reg_2[872]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1743]),.i2(intermediate_reg_1[1742]),.o(intermediate_reg_2[871]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1741]),.i2(intermediate_reg_1[1740]),.o(intermediate_reg_2[870]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1739]),.i2(intermediate_reg_1[1738]),.o(intermediate_reg_2[869]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1737]),.i2(intermediate_reg_1[1736]),.o(intermediate_reg_2[868])); 
mux_module mux_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1735]),.i2(intermediate_reg_1[1734]),.o(intermediate_reg_2[867]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1733]),.i2(intermediate_reg_1[1732]),.o(intermediate_reg_2[866]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1731]),.i2(intermediate_reg_1[1730]),.o(intermediate_reg_2[865])); 
mux_module mux_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1729]),.i2(intermediate_reg_1[1728]),.o(intermediate_reg_2[864]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1727]),.i2(intermediate_reg_1[1726]),.o(intermediate_reg_2[863])); 
mux_module mux_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1725]),.i2(intermediate_reg_1[1724]),.o(intermediate_reg_2[862]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1723]),.i2(intermediate_reg_1[1722]),.o(intermediate_reg_2[861])); 
mux_module mux_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1721]),.i2(intermediate_reg_1[1720]),.o(intermediate_reg_2[860]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1719]),.i2(intermediate_reg_1[1718]),.o(intermediate_reg_2[859])); 
mux_module mux_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1717]),.i2(intermediate_reg_1[1716]),.o(intermediate_reg_2[858]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1715]),.i2(intermediate_reg_1[1714]),.o(intermediate_reg_2[857])); 
xor_module xor_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1713]),.i2(intermediate_reg_1[1712]),.o(intermediate_reg_2[856])); 
xor_module xor_module_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1711]),.i2(intermediate_reg_1[1710]),.o(intermediate_reg_2[855])); 
mux_module mux_module_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1709]),.i2(intermediate_reg_1[1708]),.o(intermediate_reg_2[854]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1707]),.i2(intermediate_reg_1[1706]),.o(intermediate_reg_2[853]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1705]),.i2(intermediate_reg_1[1704]),.o(intermediate_reg_2[852])); 
xor_module xor_module_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1703]),.i2(intermediate_reg_1[1702]),.o(intermediate_reg_2[851])); 
xor_module xor_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1701]),.i2(intermediate_reg_1[1700]),.o(intermediate_reg_2[850])); 
mux_module mux_module_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1699]),.i2(intermediate_reg_1[1698]),.o(intermediate_reg_2[849]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1697]),.i2(intermediate_reg_1[1696]),.o(intermediate_reg_2[848])); 
xor_module xor_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1695]),.i2(intermediate_reg_1[1694]),.o(intermediate_reg_2[847])); 
xor_module xor_module_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1693]),.i2(intermediate_reg_1[1692]),.o(intermediate_reg_2[846])); 
xor_module xor_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1691]),.i2(intermediate_reg_1[1690]),.o(intermediate_reg_2[845])); 
xor_module xor_module_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1689]),.i2(intermediate_reg_1[1688]),.o(intermediate_reg_2[844])); 
xor_module xor_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1687]),.i2(intermediate_reg_1[1686]),.o(intermediate_reg_2[843])); 
xor_module xor_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1685]),.i2(intermediate_reg_1[1684]),.o(intermediate_reg_2[842])); 
xor_module xor_module_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1683]),.i2(intermediate_reg_1[1682]),.o(intermediate_reg_2[841])); 
xor_module xor_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1681]),.i2(intermediate_reg_1[1680]),.o(intermediate_reg_2[840])); 
mux_module mux_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1679]),.i2(intermediate_reg_1[1678]),.o(intermediate_reg_2[839]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1677]),.i2(intermediate_reg_1[1676]),.o(intermediate_reg_2[838]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1675]),.i2(intermediate_reg_1[1674]),.o(intermediate_reg_2[837]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1673]),.i2(intermediate_reg_1[1672]),.o(intermediate_reg_2[836]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1671]),.i2(intermediate_reg_1[1670]),.o(intermediate_reg_2[835]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1669]),.i2(intermediate_reg_1[1668]),.o(intermediate_reg_2[834])); 
mux_module mux_module_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1667]),.i2(intermediate_reg_1[1666]),.o(intermediate_reg_2[833]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1665]),.i2(intermediate_reg_1[1664]),.o(intermediate_reg_2[832]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1663]),.i2(intermediate_reg_1[1662]),.o(intermediate_reg_2[831]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1661]),.i2(intermediate_reg_1[1660]),.o(intermediate_reg_2[830]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1659]),.i2(intermediate_reg_1[1658]),.o(intermediate_reg_2[829]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1657]),.i2(intermediate_reg_1[1656]),.o(intermediate_reg_2[828]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1655]),.i2(intermediate_reg_1[1654]),.o(intermediate_reg_2[827]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1653]),.i2(intermediate_reg_1[1652]),.o(intermediate_reg_2[826]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1651]),.i2(intermediate_reg_1[1650]),.o(intermediate_reg_2[825])); 
mux_module mux_module_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1649]),.i2(intermediate_reg_1[1648]),.o(intermediate_reg_2[824]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1647]),.i2(intermediate_reg_1[1646]),.o(intermediate_reg_2[823])); 
xor_module xor_module_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1645]),.i2(intermediate_reg_1[1644]),.o(intermediate_reg_2[822])); 
mux_module mux_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1643]),.i2(intermediate_reg_1[1642]),.o(intermediate_reg_2[821]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1641]),.i2(intermediate_reg_1[1640]),.o(intermediate_reg_2[820])); 
mux_module mux_module_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1639]),.i2(intermediate_reg_1[1638]),.o(intermediate_reg_2[819]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1637]),.i2(intermediate_reg_1[1636]),.o(intermediate_reg_2[818]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1635]),.i2(intermediate_reg_1[1634]),.o(intermediate_reg_2[817])); 
mux_module mux_module_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1633]),.i2(intermediate_reg_1[1632]),.o(intermediate_reg_2[816]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1631]),.i2(intermediate_reg_1[1630]),.o(intermediate_reg_2[815]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1629]),.i2(intermediate_reg_1[1628]),.o(intermediate_reg_2[814]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1627]),.i2(intermediate_reg_1[1626]),.o(intermediate_reg_2[813]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1625]),.i2(intermediate_reg_1[1624]),.o(intermediate_reg_2[812])); 
xor_module xor_module_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1623]),.i2(intermediate_reg_1[1622]),.o(intermediate_reg_2[811])); 
xor_module xor_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1621]),.i2(intermediate_reg_1[1620]),.o(intermediate_reg_2[810])); 
mux_module mux_module_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1619]),.i2(intermediate_reg_1[1618]),.o(intermediate_reg_2[809]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1617]),.i2(intermediate_reg_1[1616]),.o(intermediate_reg_2[808]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1615]),.i2(intermediate_reg_1[1614]),.o(intermediate_reg_2[807]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1613]),.i2(intermediate_reg_1[1612]),.o(intermediate_reg_2[806]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1611]),.i2(intermediate_reg_1[1610]),.o(intermediate_reg_2[805])); 
xor_module xor_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1609]),.i2(intermediate_reg_1[1608]),.o(intermediate_reg_2[804])); 
mux_module mux_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1607]),.i2(intermediate_reg_1[1606]),.o(intermediate_reg_2[803]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1605]),.i2(intermediate_reg_1[1604]),.o(intermediate_reg_2[802]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1603]),.i2(intermediate_reg_1[1602]),.o(intermediate_reg_2[801]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1601]),.i2(intermediate_reg_1[1600]),.o(intermediate_reg_2[800]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1599]),.i2(intermediate_reg_1[1598]),.o(intermediate_reg_2[799]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1597]),.i2(intermediate_reg_1[1596]),.o(intermediate_reg_2[798]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1595]),.i2(intermediate_reg_1[1594]),.o(intermediate_reg_2[797]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1593]),.i2(intermediate_reg_1[1592]),.o(intermediate_reg_2[796]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1591]),.i2(intermediate_reg_1[1590]),.o(intermediate_reg_2[795]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1589]),.i2(intermediate_reg_1[1588]),.o(intermediate_reg_2[794])); 
mux_module mux_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1587]),.i2(intermediate_reg_1[1586]),.o(intermediate_reg_2[793]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1585]),.i2(intermediate_reg_1[1584]),.o(intermediate_reg_2[792])); 
mux_module mux_module_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1583]),.i2(intermediate_reg_1[1582]),.o(intermediate_reg_2[791]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1581]),.i2(intermediate_reg_1[1580]),.o(intermediate_reg_2[790]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1579]),.i2(intermediate_reg_1[1578]),.o(intermediate_reg_2[789])); 
mux_module mux_module_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1577]),.i2(intermediate_reg_1[1576]),.o(intermediate_reg_2[788]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1575]),.i2(intermediate_reg_1[1574]),.o(intermediate_reg_2[787]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1573]),.i2(intermediate_reg_1[1572]),.o(intermediate_reg_2[786])); 
xor_module xor_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1571]),.i2(intermediate_reg_1[1570]),.o(intermediate_reg_2[785])); 
xor_module xor_module_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1569]),.i2(intermediate_reg_1[1568]),.o(intermediate_reg_2[784])); 
xor_module xor_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1567]),.i2(intermediate_reg_1[1566]),.o(intermediate_reg_2[783])); 
xor_module xor_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1565]),.i2(intermediate_reg_1[1564]),.o(intermediate_reg_2[782])); 
xor_module xor_module_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1563]),.i2(intermediate_reg_1[1562]),.o(intermediate_reg_2[781])); 
xor_module xor_module_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1561]),.i2(intermediate_reg_1[1560]),.o(intermediate_reg_2[780])); 
mux_module mux_module_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1559]),.i2(intermediate_reg_1[1558]),.o(intermediate_reg_2[779]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1557]),.i2(intermediate_reg_1[1556]),.o(intermediate_reg_2[778])); 
xor_module xor_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1555]),.i2(intermediate_reg_1[1554]),.o(intermediate_reg_2[777])); 
mux_module mux_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1553]),.i2(intermediate_reg_1[1552]),.o(intermediate_reg_2[776]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1551]),.i2(intermediate_reg_1[1550]),.o(intermediate_reg_2[775])); 
mux_module mux_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1549]),.i2(intermediate_reg_1[1548]),.o(intermediate_reg_2[774]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1547]),.i2(intermediate_reg_1[1546]),.o(intermediate_reg_2[773]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1545]),.i2(intermediate_reg_1[1544]),.o(intermediate_reg_2[772]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1543]),.i2(intermediate_reg_1[1542]),.o(intermediate_reg_2[771]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1541]),.i2(intermediate_reg_1[1540]),.o(intermediate_reg_2[770]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1539]),.i2(intermediate_reg_1[1538]),.o(intermediate_reg_2[769]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1537]),.i2(intermediate_reg_1[1536]),.o(intermediate_reg_2[768])); 
xor_module xor_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1535]),.i2(intermediate_reg_1[1534]),.o(intermediate_reg_2[767])); 
xor_module xor_module_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1533]),.i2(intermediate_reg_1[1532]),.o(intermediate_reg_2[766])); 
mux_module mux_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1531]),.i2(intermediate_reg_1[1530]),.o(intermediate_reg_2[765]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1529]),.i2(intermediate_reg_1[1528]),.o(intermediate_reg_2[764]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1527]),.i2(intermediate_reg_1[1526]),.o(intermediate_reg_2[763])); 
mux_module mux_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1525]),.i2(intermediate_reg_1[1524]),.o(intermediate_reg_2[762]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1523]),.i2(intermediate_reg_1[1522]),.o(intermediate_reg_2[761])); 
mux_module mux_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1521]),.i2(intermediate_reg_1[1520]),.o(intermediate_reg_2[760]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1519]),.i2(intermediate_reg_1[1518]),.o(intermediate_reg_2[759]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1517]),.i2(intermediate_reg_1[1516]),.o(intermediate_reg_2[758])); 
xor_module xor_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1515]),.i2(intermediate_reg_1[1514]),.o(intermediate_reg_2[757])); 
mux_module mux_module_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1513]),.i2(intermediate_reg_1[1512]),.o(intermediate_reg_2[756]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1511]),.i2(intermediate_reg_1[1510]),.o(intermediate_reg_2[755])); 
xor_module xor_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1509]),.i2(intermediate_reg_1[1508]),.o(intermediate_reg_2[754])); 
mux_module mux_module_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1507]),.i2(intermediate_reg_1[1506]),.o(intermediate_reg_2[753]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1505]),.i2(intermediate_reg_1[1504]),.o(intermediate_reg_2[752]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1503]),.i2(intermediate_reg_1[1502]),.o(intermediate_reg_2[751]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1501]),.i2(intermediate_reg_1[1500]),.o(intermediate_reg_2[750])); 
xor_module xor_module_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1499]),.i2(intermediate_reg_1[1498]),.o(intermediate_reg_2[749])); 
mux_module mux_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1497]),.i2(intermediate_reg_1[1496]),.o(intermediate_reg_2[748]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1495]),.i2(intermediate_reg_1[1494]),.o(intermediate_reg_2[747])); 
xor_module xor_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1493]),.i2(intermediate_reg_1[1492]),.o(intermediate_reg_2[746])); 
mux_module mux_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1491]),.i2(intermediate_reg_1[1490]),.o(intermediate_reg_2[745]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1489]),.i2(intermediate_reg_1[1488]),.o(intermediate_reg_2[744])); 
mux_module mux_module_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1487]),.i2(intermediate_reg_1[1486]),.o(intermediate_reg_2[743]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1485]),.i2(intermediate_reg_1[1484]),.o(intermediate_reg_2[742]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1483]),.i2(intermediate_reg_1[1482]),.o(intermediate_reg_2[741]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1481]),.i2(intermediate_reg_1[1480]),.o(intermediate_reg_2[740]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1479]),.i2(intermediate_reg_1[1478]),.o(intermediate_reg_2[739])); 
xor_module xor_module_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1477]),.i2(intermediate_reg_1[1476]),.o(intermediate_reg_2[738])); 
mux_module mux_module_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1475]),.i2(intermediate_reg_1[1474]),.o(intermediate_reg_2[737]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1473]),.i2(intermediate_reg_1[1472]),.o(intermediate_reg_2[736])); 
mux_module mux_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1471]),.i2(intermediate_reg_1[1470]),.o(intermediate_reg_2[735]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1469]),.i2(intermediate_reg_1[1468]),.o(intermediate_reg_2[734]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1467]),.i2(intermediate_reg_1[1466]),.o(intermediate_reg_2[733])); 
xor_module xor_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1465]),.i2(intermediate_reg_1[1464]),.o(intermediate_reg_2[732])); 
mux_module mux_module_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1463]),.i2(intermediate_reg_1[1462]),.o(intermediate_reg_2[731]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1461]),.i2(intermediate_reg_1[1460]),.o(intermediate_reg_2[730]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1459]),.i2(intermediate_reg_1[1458]),.o(intermediate_reg_2[729])); 
xor_module xor_module_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1457]),.i2(intermediate_reg_1[1456]),.o(intermediate_reg_2[728])); 
mux_module mux_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1455]),.i2(intermediate_reg_1[1454]),.o(intermediate_reg_2[727]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1453]),.i2(intermediate_reg_1[1452]),.o(intermediate_reg_2[726]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1451]),.i2(intermediate_reg_1[1450]),.o(intermediate_reg_2[725]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1449]),.i2(intermediate_reg_1[1448]),.o(intermediate_reg_2[724]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1447]),.i2(intermediate_reg_1[1446]),.o(intermediate_reg_2[723])); 
xor_module xor_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1445]),.i2(intermediate_reg_1[1444]),.o(intermediate_reg_2[722])); 
xor_module xor_module_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1443]),.i2(intermediate_reg_1[1442]),.o(intermediate_reg_2[721])); 
xor_module xor_module_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1441]),.i2(intermediate_reg_1[1440]),.o(intermediate_reg_2[720])); 
xor_module xor_module_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1439]),.i2(intermediate_reg_1[1438]),.o(intermediate_reg_2[719])); 
xor_module xor_module_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1437]),.i2(intermediate_reg_1[1436]),.o(intermediate_reg_2[718])); 
xor_module xor_module_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1435]),.i2(intermediate_reg_1[1434]),.o(intermediate_reg_2[717])); 
mux_module mux_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1433]),.i2(intermediate_reg_1[1432]),.o(intermediate_reg_2[716]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1431]),.i2(intermediate_reg_1[1430]),.o(intermediate_reg_2[715])); 
xor_module xor_module_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1429]),.i2(intermediate_reg_1[1428]),.o(intermediate_reg_2[714])); 
mux_module mux_module_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1427]),.i2(intermediate_reg_1[1426]),.o(intermediate_reg_2[713]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1425]),.i2(intermediate_reg_1[1424]),.o(intermediate_reg_2[712])); 
xor_module xor_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1423]),.i2(intermediate_reg_1[1422]),.o(intermediate_reg_2[711])); 
xor_module xor_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1421]),.i2(intermediate_reg_1[1420]),.o(intermediate_reg_2[710])); 
xor_module xor_module_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1419]),.i2(intermediate_reg_1[1418]),.o(intermediate_reg_2[709])); 
xor_module xor_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1417]),.i2(intermediate_reg_1[1416]),.o(intermediate_reg_2[708])); 
xor_module xor_module_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1415]),.i2(intermediate_reg_1[1414]),.o(intermediate_reg_2[707])); 
xor_module xor_module_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1413]),.i2(intermediate_reg_1[1412]),.o(intermediate_reg_2[706])); 
xor_module xor_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1411]),.i2(intermediate_reg_1[1410]),.o(intermediate_reg_2[705])); 
xor_module xor_module_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1409]),.i2(intermediate_reg_1[1408]),.o(intermediate_reg_2[704])); 
xor_module xor_module_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1407]),.i2(intermediate_reg_1[1406]),.o(intermediate_reg_2[703])); 
mux_module mux_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1405]),.i2(intermediate_reg_1[1404]),.o(intermediate_reg_2[702]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1403]),.i2(intermediate_reg_1[1402]),.o(intermediate_reg_2[701]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1401]),.i2(intermediate_reg_1[1400]),.o(intermediate_reg_2[700])); 
mux_module mux_module_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1399]),.i2(intermediate_reg_1[1398]),.o(intermediate_reg_2[699]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1397]),.i2(intermediate_reg_1[1396]),.o(intermediate_reg_2[698]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1395]),.i2(intermediate_reg_1[1394]),.o(intermediate_reg_2[697])); 
mux_module mux_module_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1393]),.i2(intermediate_reg_1[1392]),.o(intermediate_reg_2[696]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1391]),.i2(intermediate_reg_1[1390]),.o(intermediate_reg_2[695])); 
mux_module mux_module_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1389]),.i2(intermediate_reg_1[1388]),.o(intermediate_reg_2[694]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1387]),.i2(intermediate_reg_1[1386]),.o(intermediate_reg_2[693])); 
xor_module xor_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1385]),.i2(intermediate_reg_1[1384]),.o(intermediate_reg_2[692])); 
xor_module xor_module_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1383]),.i2(intermediate_reg_1[1382]),.o(intermediate_reg_2[691])); 
mux_module mux_module_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1381]),.i2(intermediate_reg_1[1380]),.o(intermediate_reg_2[690]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1379]),.i2(intermediate_reg_1[1378]),.o(intermediate_reg_2[689]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1377]),.i2(intermediate_reg_1[1376]),.o(intermediate_reg_2[688]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1375]),.i2(intermediate_reg_1[1374]),.o(intermediate_reg_2[687])); 
xor_module xor_module_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1373]),.i2(intermediate_reg_1[1372]),.o(intermediate_reg_2[686])); 
xor_module xor_module_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1371]),.i2(intermediate_reg_1[1370]),.o(intermediate_reg_2[685])); 
xor_module xor_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1369]),.i2(intermediate_reg_1[1368]),.o(intermediate_reg_2[684])); 
xor_module xor_module_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1367]),.i2(intermediate_reg_1[1366]),.o(intermediate_reg_2[683])); 
xor_module xor_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1365]),.i2(intermediate_reg_1[1364]),.o(intermediate_reg_2[682])); 
xor_module xor_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1363]),.i2(intermediate_reg_1[1362]),.o(intermediate_reg_2[681])); 
xor_module xor_module_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1361]),.i2(intermediate_reg_1[1360]),.o(intermediate_reg_2[680])); 
xor_module xor_module_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1359]),.i2(intermediate_reg_1[1358]),.o(intermediate_reg_2[679])); 
xor_module xor_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1357]),.i2(intermediate_reg_1[1356]),.o(intermediate_reg_2[678])); 
mux_module mux_module_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1355]),.i2(intermediate_reg_1[1354]),.o(intermediate_reg_2[677]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1353]),.i2(intermediate_reg_1[1352]),.o(intermediate_reg_2[676])); 
mux_module mux_module_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1351]),.i2(intermediate_reg_1[1350]),.o(intermediate_reg_2[675]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1349]),.i2(intermediate_reg_1[1348]),.o(intermediate_reg_2[674])); 
mux_module mux_module_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1347]),.i2(intermediate_reg_1[1346]),.o(intermediate_reg_2[673]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1345]),.i2(intermediate_reg_1[1344]),.o(intermediate_reg_2[672])); 
mux_module mux_module_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1343]),.i2(intermediate_reg_1[1342]),.o(intermediate_reg_2[671]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1341]),.i2(intermediate_reg_1[1340]),.o(intermediate_reg_2[670])); 
mux_module mux_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1339]),.i2(intermediate_reg_1[1338]),.o(intermediate_reg_2[669]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1337]),.i2(intermediate_reg_1[1336]),.o(intermediate_reg_2[668])); 
xor_module xor_module_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1335]),.i2(intermediate_reg_1[1334]),.o(intermediate_reg_2[667])); 
xor_module xor_module_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1333]),.i2(intermediate_reg_1[1332]),.o(intermediate_reg_2[666])); 
mux_module mux_module_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1331]),.i2(intermediate_reg_1[1330]),.o(intermediate_reg_2[665]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1329]),.i2(intermediate_reg_1[1328]),.o(intermediate_reg_2[664]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1327]),.i2(intermediate_reg_1[1326]),.o(intermediate_reg_2[663])); 
mux_module mux_module_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1325]),.i2(intermediate_reg_1[1324]),.o(intermediate_reg_2[662]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1323]),.i2(intermediate_reg_1[1322]),.o(intermediate_reg_2[661]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1321]),.i2(intermediate_reg_1[1320]),.o(intermediate_reg_2[660])); 
xor_module xor_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1319]),.i2(intermediate_reg_1[1318]),.o(intermediate_reg_2[659])); 
mux_module mux_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1317]),.i2(intermediate_reg_1[1316]),.o(intermediate_reg_2[658]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1315]),.i2(intermediate_reg_1[1314]),.o(intermediate_reg_2[657]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1313]),.i2(intermediate_reg_1[1312]),.o(intermediate_reg_2[656])); 
xor_module xor_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1311]),.i2(intermediate_reg_1[1310]),.o(intermediate_reg_2[655])); 
xor_module xor_module_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1309]),.i2(intermediate_reg_1[1308]),.o(intermediate_reg_2[654])); 
mux_module mux_module_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1307]),.i2(intermediate_reg_1[1306]),.o(intermediate_reg_2[653]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1305]),.i2(intermediate_reg_1[1304]),.o(intermediate_reg_2[652]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1303]),.i2(intermediate_reg_1[1302]),.o(intermediate_reg_2[651])); 
xor_module xor_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1301]),.i2(intermediate_reg_1[1300]),.o(intermediate_reg_2[650])); 
mux_module mux_module_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1299]),.i2(intermediate_reg_1[1298]),.o(intermediate_reg_2[649]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1297]),.i2(intermediate_reg_1[1296]),.o(intermediate_reg_2[648])); 
xor_module xor_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1295]),.i2(intermediate_reg_1[1294]),.o(intermediate_reg_2[647])); 
mux_module mux_module_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1293]),.i2(intermediate_reg_1[1292]),.o(intermediate_reg_2[646]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1291]),.i2(intermediate_reg_1[1290]),.o(intermediate_reg_2[645]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1289]),.i2(intermediate_reg_1[1288]),.o(intermediate_reg_2[644])); 
mux_module mux_module_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1287]),.i2(intermediate_reg_1[1286]),.o(intermediate_reg_2[643]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1285]),.i2(intermediate_reg_1[1284]),.o(intermediate_reg_2[642])); 
mux_module mux_module_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1283]),.i2(intermediate_reg_1[1282]),.o(intermediate_reg_2[641]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1281]),.i2(intermediate_reg_1[1280]),.o(intermediate_reg_2[640])); 
mux_module mux_module_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1279]),.i2(intermediate_reg_1[1278]),.o(intermediate_reg_2[639]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1277]),.i2(intermediate_reg_1[1276]),.o(intermediate_reg_2[638])); 
xor_module xor_module_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1275]),.i2(intermediate_reg_1[1274]),.o(intermediate_reg_2[637])); 
xor_module xor_module_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1273]),.i2(intermediate_reg_1[1272]),.o(intermediate_reg_2[636])); 
xor_module xor_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1271]),.i2(intermediate_reg_1[1270]),.o(intermediate_reg_2[635])); 
mux_module mux_module_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1269]),.i2(intermediate_reg_1[1268]),.o(intermediate_reg_2[634]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1267]),.i2(intermediate_reg_1[1266]),.o(intermediate_reg_2[633])); 
xor_module xor_module_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1265]),.i2(intermediate_reg_1[1264]),.o(intermediate_reg_2[632])); 
xor_module xor_module_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1263]),.i2(intermediate_reg_1[1262]),.o(intermediate_reg_2[631])); 
xor_module xor_module_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1261]),.i2(intermediate_reg_1[1260]),.o(intermediate_reg_2[630])); 
xor_module xor_module_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1259]),.i2(intermediate_reg_1[1258]),.o(intermediate_reg_2[629])); 
mux_module mux_module_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1257]),.i2(intermediate_reg_1[1256]),.o(intermediate_reg_2[628]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1255]),.i2(intermediate_reg_1[1254]),.o(intermediate_reg_2[627]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1253]),.i2(intermediate_reg_1[1252]),.o(intermediate_reg_2[626]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1251]),.i2(intermediate_reg_1[1250]),.o(intermediate_reg_2[625])); 
mux_module mux_module_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1249]),.i2(intermediate_reg_1[1248]),.o(intermediate_reg_2[624]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1247]),.i2(intermediate_reg_1[1246]),.o(intermediate_reg_2[623])); 
xor_module xor_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1245]),.i2(intermediate_reg_1[1244]),.o(intermediate_reg_2[622])); 
xor_module xor_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1243]),.i2(intermediate_reg_1[1242]),.o(intermediate_reg_2[621])); 
xor_module xor_module_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1241]),.i2(intermediate_reg_1[1240]),.o(intermediate_reg_2[620])); 
xor_module xor_module_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1239]),.i2(intermediate_reg_1[1238]),.o(intermediate_reg_2[619])); 
xor_module xor_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1237]),.i2(intermediate_reg_1[1236]),.o(intermediate_reg_2[618])); 
mux_module mux_module_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1235]),.i2(intermediate_reg_1[1234]),.o(intermediate_reg_2[617]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1233]),.i2(intermediate_reg_1[1232]),.o(intermediate_reg_2[616])); 
xor_module xor_module_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1231]),.i2(intermediate_reg_1[1230]),.o(intermediate_reg_2[615])); 
xor_module xor_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1229]),.i2(intermediate_reg_1[1228]),.o(intermediate_reg_2[614])); 
xor_module xor_module_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1227]),.i2(intermediate_reg_1[1226]),.o(intermediate_reg_2[613])); 
mux_module mux_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1225]),.i2(intermediate_reg_1[1224]),.o(intermediate_reg_2[612]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1223]),.i2(intermediate_reg_1[1222]),.o(intermediate_reg_2[611])); 
xor_module xor_module_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1221]),.i2(intermediate_reg_1[1220]),.o(intermediate_reg_2[610])); 
mux_module mux_module_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1219]),.i2(intermediate_reg_1[1218]),.o(intermediate_reg_2[609]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1217]),.i2(intermediate_reg_1[1216]),.o(intermediate_reg_2[608]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1215]),.i2(intermediate_reg_1[1214]),.o(intermediate_reg_2[607]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1213]),.i2(intermediate_reg_1[1212]),.o(intermediate_reg_2[606]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1211]),.i2(intermediate_reg_1[1210]),.o(intermediate_reg_2[605]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1209]),.i2(intermediate_reg_1[1208]),.o(intermediate_reg_2[604])); 
xor_module xor_module_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1207]),.i2(intermediate_reg_1[1206]),.o(intermediate_reg_2[603])); 
xor_module xor_module_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1205]),.i2(intermediate_reg_1[1204]),.o(intermediate_reg_2[602])); 
xor_module xor_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1203]),.i2(intermediate_reg_1[1202]),.o(intermediate_reg_2[601])); 
mux_module mux_module_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1201]),.i2(intermediate_reg_1[1200]),.o(intermediate_reg_2[600]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1199]),.i2(intermediate_reg_1[1198]),.o(intermediate_reg_2[599])); 
xor_module xor_module_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1197]),.i2(intermediate_reg_1[1196]),.o(intermediate_reg_2[598])); 
xor_module xor_module_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1195]),.i2(intermediate_reg_1[1194]),.o(intermediate_reg_2[597])); 
xor_module xor_module_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1193]),.i2(intermediate_reg_1[1192]),.o(intermediate_reg_2[596])); 
xor_module xor_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1191]),.i2(intermediate_reg_1[1190]),.o(intermediate_reg_2[595])); 
mux_module mux_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1189]),.i2(intermediate_reg_1[1188]),.o(intermediate_reg_2[594]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1187]),.i2(intermediate_reg_1[1186]),.o(intermediate_reg_2[593])); 
mux_module mux_module_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1185]),.i2(intermediate_reg_1[1184]),.o(intermediate_reg_2[592]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1183]),.i2(intermediate_reg_1[1182]),.o(intermediate_reg_2[591]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1181]),.i2(intermediate_reg_1[1180]),.o(intermediate_reg_2[590])); 
mux_module mux_module_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1179]),.i2(intermediate_reg_1[1178]),.o(intermediate_reg_2[589]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1177]),.i2(intermediate_reg_1[1176]),.o(intermediate_reg_2[588]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1175]),.i2(intermediate_reg_1[1174]),.o(intermediate_reg_2[587]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1173]),.i2(intermediate_reg_1[1172]),.o(intermediate_reg_2[586])); 
mux_module mux_module_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1171]),.i2(intermediate_reg_1[1170]),.o(intermediate_reg_2[585]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1169]),.i2(intermediate_reg_1[1168]),.o(intermediate_reg_2[584])); 
mux_module mux_module_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1167]),.i2(intermediate_reg_1[1166]),.o(intermediate_reg_2[583]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1165]),.i2(intermediate_reg_1[1164]),.o(intermediate_reg_2[582]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1163]),.i2(intermediate_reg_1[1162]),.o(intermediate_reg_2[581])); 
mux_module mux_module_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1161]),.i2(intermediate_reg_1[1160]),.o(intermediate_reg_2[580]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1159]),.i2(intermediate_reg_1[1158]),.o(intermediate_reg_2[579]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1157]),.i2(intermediate_reg_1[1156]),.o(intermediate_reg_2[578]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1155]),.i2(intermediate_reg_1[1154]),.o(intermediate_reg_2[577]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1153]),.i2(intermediate_reg_1[1152]),.o(intermediate_reg_2[576]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1151]),.i2(intermediate_reg_1[1150]),.o(intermediate_reg_2[575])); 
xor_module xor_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1149]),.i2(intermediate_reg_1[1148]),.o(intermediate_reg_2[574])); 
xor_module xor_module_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1147]),.i2(intermediate_reg_1[1146]),.o(intermediate_reg_2[573])); 
mux_module mux_module_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1145]),.i2(intermediate_reg_1[1144]),.o(intermediate_reg_2[572]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1143]),.i2(intermediate_reg_1[1142]),.o(intermediate_reg_2[571])); 
xor_module xor_module_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1141]),.i2(intermediate_reg_1[1140]),.o(intermediate_reg_2[570])); 
xor_module xor_module_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1139]),.i2(intermediate_reg_1[1138]),.o(intermediate_reg_2[569])); 
mux_module mux_module_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1137]),.i2(intermediate_reg_1[1136]),.o(intermediate_reg_2[568]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1135]),.i2(intermediate_reg_1[1134]),.o(intermediate_reg_2[567]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1133]),.i2(intermediate_reg_1[1132]),.o(intermediate_reg_2[566])); 
mux_module mux_module_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1131]),.i2(intermediate_reg_1[1130]),.o(intermediate_reg_2[565]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1129]),.i2(intermediate_reg_1[1128]),.o(intermediate_reg_2[564])); 
mux_module mux_module_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1127]),.i2(intermediate_reg_1[1126]),.o(intermediate_reg_2[563]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1125]),.i2(intermediate_reg_1[1124]),.o(intermediate_reg_2[562]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1123]),.i2(intermediate_reg_1[1122]),.o(intermediate_reg_2[561])); 
xor_module xor_module_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1121]),.i2(intermediate_reg_1[1120]),.o(intermediate_reg_2[560])); 
mux_module mux_module_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1119]),.i2(intermediate_reg_1[1118]),.o(intermediate_reg_2[559]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1117]),.i2(intermediate_reg_1[1116]),.o(intermediate_reg_2[558])); 
mux_module mux_module_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1115]),.i2(intermediate_reg_1[1114]),.o(intermediate_reg_2[557]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1113]),.i2(intermediate_reg_1[1112]),.o(intermediate_reg_2[556])); 
xor_module xor_module_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1111]),.i2(intermediate_reg_1[1110]),.o(intermediate_reg_2[555])); 
mux_module mux_module_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1109]),.i2(intermediate_reg_1[1108]),.o(intermediate_reg_2[554]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1107]),.i2(intermediate_reg_1[1106]),.o(intermediate_reg_2[553])); 
mux_module mux_module_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1105]),.i2(intermediate_reg_1[1104]),.o(intermediate_reg_2[552]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1103]),.i2(intermediate_reg_1[1102]),.o(intermediate_reg_2[551]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1101]),.i2(intermediate_reg_1[1100]),.o(intermediate_reg_2[550]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1099]),.i2(intermediate_reg_1[1098]),.o(intermediate_reg_2[549]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1097]),.i2(intermediate_reg_1[1096]),.o(intermediate_reg_2[548]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1095]),.i2(intermediate_reg_1[1094]),.o(intermediate_reg_2[547])); 
xor_module xor_module_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1093]),.i2(intermediate_reg_1[1092]),.o(intermediate_reg_2[546])); 
mux_module mux_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1091]),.i2(intermediate_reg_1[1090]),.o(intermediate_reg_2[545]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1089]),.i2(intermediate_reg_1[1088]),.o(intermediate_reg_2[544]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1087]),.i2(intermediate_reg_1[1086]),.o(intermediate_reg_2[543]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1085]),.i2(intermediate_reg_1[1084]),.o(intermediate_reg_2[542])); 
mux_module mux_module_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1083]),.i2(intermediate_reg_1[1082]),.o(intermediate_reg_2[541]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1081]),.i2(intermediate_reg_1[1080]),.o(intermediate_reg_2[540]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1079]),.i2(intermediate_reg_1[1078]),.o(intermediate_reg_2[539])); 
mux_module mux_module_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1077]),.i2(intermediate_reg_1[1076]),.o(intermediate_reg_2[538]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1075]),.i2(intermediate_reg_1[1074]),.o(intermediate_reg_2[537]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1073]),.i2(intermediate_reg_1[1072]),.o(intermediate_reg_2[536]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1071]),.i2(intermediate_reg_1[1070]),.o(intermediate_reg_2[535]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1069]),.i2(intermediate_reg_1[1068]),.o(intermediate_reg_2[534]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1067]),.i2(intermediate_reg_1[1066]),.o(intermediate_reg_2[533])); 
mux_module mux_module_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1065]),.i2(intermediate_reg_1[1064]),.o(intermediate_reg_2[532]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1063]),.i2(intermediate_reg_1[1062]),.o(intermediate_reg_2[531])); 
xor_module xor_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1061]),.i2(intermediate_reg_1[1060]),.o(intermediate_reg_2[530])); 
mux_module mux_module_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1059]),.i2(intermediate_reg_1[1058]),.o(intermediate_reg_2[529]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1057]),.i2(intermediate_reg_1[1056]),.o(intermediate_reg_2[528])); 
xor_module xor_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1055]),.i2(intermediate_reg_1[1054]),.o(intermediate_reg_2[527])); 
mux_module mux_module_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1053]),.i2(intermediate_reg_1[1052]),.o(intermediate_reg_2[526]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1051]),.i2(intermediate_reg_1[1050]),.o(intermediate_reg_2[525]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1049]),.i2(intermediate_reg_1[1048]),.o(intermediate_reg_2[524]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1047]),.i2(intermediate_reg_1[1046]),.o(intermediate_reg_2[523])); 
xor_module xor_module_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1045]),.i2(intermediate_reg_1[1044]),.o(intermediate_reg_2[522])); 
mux_module mux_module_inst_2_514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1043]),.i2(intermediate_reg_1[1042]),.o(intermediate_reg_2[521]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1041]),.i2(intermediate_reg_1[1040]),.o(intermediate_reg_2[520]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1039]),.i2(intermediate_reg_1[1038]),.o(intermediate_reg_2[519])); 
mux_module mux_module_inst_2_517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1037]),.i2(intermediate_reg_1[1036]),.o(intermediate_reg_2[518]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1035]),.i2(intermediate_reg_1[1034]),.o(intermediate_reg_2[517])); 
xor_module xor_module_inst_2_519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1033]),.i2(intermediate_reg_1[1032]),.o(intermediate_reg_2[516])); 
xor_module xor_module_inst_2_520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1031]),.i2(intermediate_reg_1[1030]),.o(intermediate_reg_2[515])); 
mux_module mux_module_inst_2_521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1029]),.i2(intermediate_reg_1[1028]),.o(intermediate_reg_2[514]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512])); 
xor_module xor_module_inst_2_524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511])); 
xor_module xor_module_inst_2_525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510])); 
mux_module mux_module_inst_2_526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506])); 
mux_module mux_module_inst_2_530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504])); 
xor_module xor_module_inst_2_532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503])); 
mux_module mux_module_inst_2_533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500])); 
xor_module xor_module_inst_2_536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499])); 
mux_module mux_module_inst_2_537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497])); 
mux_module mux_module_inst_2_539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493])); 
mux_module mux_module_inst_2_543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491])); 
mux_module mux_module_inst_2_545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488])); 
xor_module xor_module_inst_2_548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487])); 
mux_module mux_module_inst_2_549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485])); 
mux_module mux_module_inst_2_551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483])); 
mux_module mux_module_inst_2_553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
mux_module mux_module_inst_2_557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_560(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_561(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_562(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473])); 
mux_module mux_module_inst_2_563(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_564(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471])); 
xor_module xor_module_inst_2_565(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470])); 
xor_module xor_module_inst_2_566(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469])); 
xor_module xor_module_inst_2_567(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468])); 
xor_module xor_module_inst_2_568(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467])); 
xor_module xor_module_inst_2_569(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466])); 
xor_module xor_module_inst_2_570(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465])); 
mux_module mux_module_inst_2_571(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_572(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_573(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_574(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_575(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460])); 
mux_module mux_module_inst_2_576(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_577(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458])); 
mux_module mux_module_inst_2_578(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_579(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456])); 
mux_module mux_module_inst_2_580(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_581(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_582(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_583(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452])); 
mux_module mux_module_inst_2_584(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_585(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450])); 
xor_module xor_module_inst_2_586(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449])); 
mux_module mux_module_inst_2_587(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_588(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447])); 
xor_module xor_module_inst_2_589(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446])); 
xor_module xor_module_inst_2_590(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445])); 
mux_module mux_module_inst_2_591(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_592(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443])); 
xor_module xor_module_inst_2_593(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442])); 
xor_module xor_module_inst_2_594(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441])); 
mux_module mux_module_inst_2_595(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_596(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_597(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_598(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437])); 
xor_module xor_module_inst_2_599(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436])); 
xor_module xor_module_inst_2_600(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435])); 
xor_module xor_module_inst_2_601(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434])); 
mux_module mux_module_inst_2_602(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_603(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432])); 
mux_module mux_module_inst_2_604(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_605(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_606(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429])); 
mux_module mux_module_inst_2_607(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_608(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427])); 
xor_module xor_module_inst_2_609(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426])); 
xor_module xor_module_inst_2_610(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425])); 
xor_module xor_module_inst_2_611(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424])); 
mux_module mux_module_inst_2_612(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_613(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_614(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421])); 
mux_module mux_module_inst_2_615(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_616(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419])); 
mux_module mux_module_inst_2_617(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_618(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_619(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416])); 
mux_module mux_module_inst_2_620(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_621(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_622(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413])); 
xor_module xor_module_inst_2_623(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412])); 
mux_module mux_module_inst_2_624(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_625(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_626(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_627(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_628(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_629(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406])); 
mux_module mux_module_inst_2_630(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_631(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404])); 
mux_module mux_module_inst_2_632(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_633(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402])); 
mux_module mux_module_inst_2_634(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_635(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_636(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_637(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_638(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397])); 
xor_module xor_module_inst_2_639(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396])); 
mux_module mux_module_inst_2_640(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_641(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_642(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_643(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392])); 
mux_module mux_module_inst_2_644(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_645(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_646(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389])); 
mux_module mux_module_inst_2_647(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_648(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387])); 
mux_module mux_module_inst_2_649(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_650(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_651(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384])); 
xor_module xor_module_inst_2_652(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383])); 
xor_module xor_module_inst_2_653(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382])); 
mux_module mux_module_inst_2_654(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_655(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
mux_module mux_module_inst_2_656(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_657(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_658(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_659(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376])); 
mux_module mux_module_inst_2_660(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_661(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_662(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_663(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_664(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_665(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
xor_module xor_module_inst_2_666(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369])); 
mux_module mux_module_inst_2_667(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_668(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367])); 
xor_module xor_module_inst_2_669(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366])); 
xor_module xor_module_inst_2_670(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365])); 
xor_module xor_module_inst_2_671(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
xor_module xor_module_inst_2_672(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363])); 
mux_module mux_module_inst_2_673(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_674(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361])); 
xor_module xor_module_inst_2_675(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360])); 
xor_module xor_module_inst_2_676(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
xor_module xor_module_inst_2_677(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
mux_module mux_module_inst_2_678(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_679(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_680(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355])); 
mux_module mux_module_inst_2_681(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_682(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353])); 
xor_module xor_module_inst_2_683(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352])); 
xor_module xor_module_inst_2_684(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351])); 
xor_module xor_module_inst_2_685(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350])); 
xor_module xor_module_inst_2_686(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349])); 
mux_module mux_module_inst_2_687(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_688(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_689(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346])); 
xor_module xor_module_inst_2_690(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345])); 
xor_module xor_module_inst_2_691(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
xor_module xor_module_inst_2_692(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343])); 
mux_module mux_module_inst_2_693(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_694(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_695(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340])); 
mux_module mux_module_inst_2_696(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_697(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338])); 
xor_module xor_module_inst_2_698(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337])); 
mux_module mux_module_inst_2_699(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_700(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_701(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334])); 
mux_module mux_module_inst_2_702(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_703(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_704(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_705(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
xor_module xor_module_inst_2_706(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
xor_module xor_module_inst_2_707(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328])); 
xor_module xor_module_inst_2_708(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
mux_module mux_module_inst_2_709(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_710(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325])); 
mux_module mux_module_inst_2_711(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_712(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323])); 
xor_module xor_module_inst_2_713(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322])); 
mux_module mux_module_inst_2_714(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_715(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
mux_module mux_module_inst_2_716(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_717(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318])); 
xor_module xor_module_inst_2_718(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317])); 
xor_module xor_module_inst_2_719(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316])); 
xor_module xor_module_inst_2_720(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315])); 
mux_module mux_module_inst_2_721(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_722(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313])); 
mux_module mux_module_inst_2_723(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_724(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_725(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_726(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_727(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308])); 
mux_module mux_module_inst_2_728(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_729(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306])); 
xor_module xor_module_inst_2_730(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305])); 
xor_module xor_module_inst_2_731(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304])); 
xor_module xor_module_inst_2_732(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
mux_module mux_module_inst_2_733(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_734(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
mux_module mux_module_inst_2_735(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_736(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_737(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_738(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_739(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
xor_module xor_module_inst_2_740(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
xor_module xor_module_inst_2_741(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294])); 
mux_module mux_module_inst_2_742(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_743(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292])); 
xor_module xor_module_inst_2_744(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291])); 
mux_module mux_module_inst_2_745(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_746(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_747(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_748(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_749(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286])); 
xor_module xor_module_inst_2_750(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
mux_module mux_module_inst_2_751(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_752(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_753(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282])); 
mux_module mux_module_inst_2_754(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_755(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280])); 
mux_module mux_module_inst_2_756(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_757(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278])); 
mux_module mux_module_inst_2_758(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_759(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276])); 
xor_module xor_module_inst_2_760(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275])); 
xor_module xor_module_inst_2_761(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
xor_module xor_module_inst_2_762(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
mux_module mux_module_inst_2_763(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_764(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_765(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270])); 
xor_module xor_module_inst_2_766(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
xor_module xor_module_inst_2_767(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268])); 
mux_module mux_module_inst_2_768(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_769(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_770(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
xor_module xor_module_inst_2_771(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264])); 
xor_module xor_module_inst_2_772(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263])); 
xor_module xor_module_inst_2_773(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
mux_module mux_module_inst_2_774(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_775(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
mux_module mux_module_inst_2_776(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_777(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_778(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_779(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
xor_module xor_module_inst_2_780(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255])); 
xor_module xor_module_inst_2_781(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254])); 
xor_module xor_module_inst_2_782(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253])); 
xor_module xor_module_inst_2_783(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252])); 
xor_module xor_module_inst_2_784(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
xor_module xor_module_inst_2_785(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250])); 
mux_module mux_module_inst_2_786(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_787(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248])); 
mux_module mux_module_inst_2_788(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_789(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246])); 
xor_module xor_module_inst_2_790(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
xor_module xor_module_inst_2_791(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244])); 
mux_module mux_module_inst_2_792(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_793(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242])); 
xor_module xor_module_inst_2_794(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
xor_module xor_module_inst_2_795(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240])); 
mux_module mux_module_inst_2_796(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_797(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
xor_module xor_module_inst_2_798(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
xor_module xor_module_inst_2_799(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236])); 
mux_module mux_module_inst_2_800(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_801(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
mux_module mux_module_inst_2_802(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_803(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_804(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231])); 
xor_module xor_module_inst_2_805(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230])); 
xor_module xor_module_inst_2_806(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229])); 
xor_module xor_module_inst_2_807(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
xor_module xor_module_inst_2_808(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227])); 
xor_module xor_module_inst_2_809(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
xor_module xor_module_inst_2_810(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
mux_module mux_module_inst_2_811(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_812(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_813(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
mux_module mux_module_inst_2_814(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_815(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_816(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_817(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
xor_module xor_module_inst_2_818(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217])); 
mux_module mux_module_inst_2_819(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_820(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215])); 
mux_module mux_module_inst_2_821(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_822(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
xor_module xor_module_inst_2_823(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
xor_module xor_module_inst_2_824(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
xor_module xor_module_inst_2_825(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
mux_module mux_module_inst_2_826(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_827(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208])); 
xor_module xor_module_inst_2_828(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
xor_module xor_module_inst_2_829(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
xor_module xor_module_inst_2_830(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
mux_module mux_module_inst_2_831(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_832(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_833(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_834(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_835(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200])); 
xor_module xor_module_inst_2_836(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
mux_module mux_module_inst_2_837(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_838(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197])); 
mux_module mux_module_inst_2_839(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_840(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_841(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_842(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193])); 
xor_module xor_module_inst_2_843(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
xor_module xor_module_inst_2_844(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
mux_module mux_module_inst_2_845(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_846(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_847(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
xor_module xor_module_inst_2_848(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
xor_module xor_module_inst_2_849(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186])); 
mux_module mux_module_inst_2_850(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_851(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
xor_module xor_module_inst_2_852(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183])); 
mux_module mux_module_inst_2_853(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_854(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_855(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180])); 
xor_module xor_module_inst_2_856(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179])); 
mux_module mux_module_inst_2_857(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_858(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
xor_module xor_module_inst_2_859(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176])); 
xor_module xor_module_inst_2_860(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175])); 
mux_module mux_module_inst_2_861(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_862(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_863(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
xor_module xor_module_inst_2_864(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
mux_module mux_module_inst_2_865(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_866(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169])); 
mux_module mux_module_inst_2_867(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_868(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167])); 
xor_module xor_module_inst_2_869(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166])); 
mux_module mux_module_inst_2_870(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_871(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_872(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
mux_module mux_module_inst_2_873(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_874(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161])); 
xor_module xor_module_inst_2_875(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160])); 
xor_module xor_module_inst_2_876(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
mux_module mux_module_inst_2_877(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_878(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_879(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156])); 
xor_module xor_module_inst_2_880(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155])); 
mux_module mux_module_inst_2_881(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_882(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_883(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_884(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_885(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
xor_module xor_module_inst_2_886(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
mux_module mux_module_inst_2_887(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_888(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147])); 
mux_module mux_module_inst_2_889(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_890(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_891(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_892(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143])); 
mux_module mux_module_inst_2_893(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_894(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_895(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_896(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_897(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138])); 
xor_module xor_module_inst_2_898(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
mux_module mux_module_inst_2_899(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_900(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135])); 
xor_module xor_module_inst_2_901(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
xor_module xor_module_inst_2_902(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133])); 
xor_module xor_module_inst_2_903(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132])); 
mux_module mux_module_inst_2_904(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_905(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130])); 
xor_module xor_module_inst_2_906(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129])); 
xor_module xor_module_inst_2_907(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
mux_module mux_module_inst_2_908(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_909(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_910(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_911(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_912(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_913(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
xor_module xor_module_inst_2_914(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121])); 
xor_module xor_module_inst_2_915(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120])); 
xor_module xor_module_inst_2_916(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119])); 
mux_module mux_module_inst_2_917(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_918(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117])); 
xor_module xor_module_inst_2_919(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116])); 
mux_module mux_module_inst_2_920(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_921(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
mux_module mux_module_inst_2_922(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_923(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
xor_module xor_module_inst_2_924(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111])); 
mux_module mux_module_inst_2_925(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_926(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_927(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
xor_module xor_module_inst_2_928(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107])); 
xor_module xor_module_inst_2_929(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
mux_module mux_module_inst_2_930(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_931(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_932(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
mux_module mux_module_inst_2_933(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_934(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_935(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100])); 
xor_module xor_module_inst_2_936(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99])); 
mux_module mux_module_inst_2_937(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_938(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
xor_module xor_module_inst_2_939(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96])); 
xor_module xor_module_inst_2_940(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95])); 
xor_module xor_module_inst_2_941(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94])); 
xor_module xor_module_inst_2_942(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
mux_module mux_module_inst_2_943(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_944(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91])); 
mux_module mux_module_inst_2_945(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_946(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_947(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_948(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_949(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
xor_module xor_module_inst_2_950(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
xor_module xor_module_inst_2_951(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
xor_module xor_module_inst_2_952(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
mux_module mux_module_inst_2_953(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_954(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
mux_module mux_module_inst_2_955(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_956(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_957(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78])); 
xor_module xor_module_inst_2_958(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
mux_module mux_module_inst_2_959(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_960(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
mux_module mux_module_inst_2_961(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_962(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73])); 
mux_module mux_module_inst_2_963(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_964(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71])); 
mux_module mux_module_inst_2_965(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_966(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69])); 
mux_module mux_module_inst_2_967(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_968(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_969(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66])); 
mux_module mux_module_inst_2_970(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_971(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_972(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
mux_module mux_module_inst_2_973(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_974(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_975(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_976(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59])); 
mux_module mux_module_inst_2_977(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_978(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_979(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56])); 
xor_module xor_module_inst_2_980(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55])); 
xor_module xor_module_inst_2_981(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54])); 
mux_module mux_module_inst_2_982(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_983(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
mux_module mux_module_inst_2_984(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_985(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
mux_module mux_module_inst_2_986(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_987(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_988(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_989(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_990(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_991(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_992(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_993(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_994(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
xor_module xor_module_inst_2_995(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40])); 
xor_module xor_module_inst_2_996(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39])); 
mux_module mux_module_inst_2_997(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_998(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_999(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35])); 
mux_module mux_module_inst_2_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33])); 
xor_module xor_module_inst_2_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32])); 
mux_module mux_module_inst_2_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
xor_module xor_module_inst_2_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29])); 
mux_module mux_module_inst_2_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27])); 
mux_module mux_module_inst_2_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22])); 
mux_module mux_module_inst_2_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20])); 
xor_module xor_module_inst_2_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
xor_module xor_module_inst_2_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18])); 
xor_module xor_module_inst_2_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17])); 
mux_module mux_module_inst_2_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14])); 
mux_module mux_module_inst_2_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
mux_module mux_module_inst_2_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5])); 
xor_module xor_module_inst_2_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
xor_module xor_module_inst_2_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
mux_module mux_module_inst_2_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
mux_module mux_module_inst_2_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0]),.sel(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [1035:0] <= intermediate_reg_2; 
outp[1319:1036] <= intermediate_reg_2[283:0] ; 
end 
endmodule 
 

module interface_14(input [2687:0] inp, output reg [1055:0] outp, input clk, input reset);
reg [2687:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1343:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342])); 
xor_module xor_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311])); 
xor_module xor_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303])); 
xor_module xor_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296])); 
mux_module mux_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292])); 
xor_module xor_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279])); 
mux_module mux_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274])); 
xor_module xor_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270])); 
xor_module xor_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262])); 
xor_module xor_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254])); 
xor_module xor_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253])); 
mux_module mux_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244])); 
mux_module mux_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
xor_module xor_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239])); 
mux_module mux_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
mux_module mux_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224])); 
xor_module xor_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
xor_module xor_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218])); 
xor_module xor_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217])); 
xor_module xor_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208])); 
xor_module xor_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206])); 
xor_module xor_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201])); 
xor_module xor_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200])); 
xor_module xor_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199])); 
xor_module xor_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197])); 
xor_module xor_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196])); 
xor_module xor_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193])); 
mux_module mux_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191])); 
mux_module mux_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186])); 
mux_module mux_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174])); 
mux_module mux_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169])); 
xor_module xor_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168])); 
mux_module mux_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165])); 
mux_module mux_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163])); 
xor_module xor_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161])); 
xor_module xor_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144])); 
xor_module xor_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141])); 
mux_module mux_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136])); 
xor_module xor_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135])); 
xor_module xor_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132])); 
mux_module mux_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
xor_module xor_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
xor_module xor_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
xor_module xor_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
xor_module xor_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118])); 
xor_module xor_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117])); 
mux_module mux_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109])); 
xor_module xor_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
mux_module mux_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
mux_module mux_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100])); 
xor_module xor_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099])); 
xor_module xor_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
xor_module xor_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084])); 
xor_module xor_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063])); 
xor_module xor_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058])); 
mux_module mux_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055])); 
xor_module xor_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
xor_module xor_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039])); 
mux_module mux_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034])); 
xor_module xor_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033])); 
xor_module xor_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
mux_module mux_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024])); 
xor_module xor_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
xor_module xor_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018])); 
xor_module xor_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
xor_module xor_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013])); 
xor_module xor_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012])); 
mux_module mux_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
xor_module xor_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999])); 
mux_module mux_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
mux_module mux_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
xor_module xor_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
mux_module mux_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
mux_module mux_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
mux_module mux_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
xor_module xor_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
mux_module mux_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
xor_module xor_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
xor_module xor_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
mux_module mux_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
xor_module xor_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
xor_module xor_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
mux_module mux_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
mux_module mux_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
xor_module xor_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
mux_module mux_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
xor_module xor_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
mux_module mux_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
xor_module xor_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
mux_module mux_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
xor_module xor_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
mux_module mux_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
xor_module xor_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
xor_module xor_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
xor_module xor_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
xor_module xor_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
xor_module xor_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
mux_module mux_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
xor_module xor_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884])); 
xor_module xor_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865])); 
xor_module xor_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
xor_module xor_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
xor_module xor_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
mux_module mux_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
xor_module xor_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
xor_module xor_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
xor_module xor_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
mux_module mux_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
mux_module mux_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842])); 
mux_module mux_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
xor_module xor_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
xor_module xor_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
xor_module xor_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
xor_module xor_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
mux_module mux_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
xor_module xor_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
xor_module xor_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
xor_module xor_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
xor_module xor_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
xor_module xor_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
xor_module xor_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
xor_module xor_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
xor_module xor_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
xor_module xor_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
xor_module xor_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
xor_module xor_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
xor_module xor_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
xor_module xor_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
xor_module xor_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
xor_module xor_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
xor_module xor_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
xor_module xor_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
mux_module mux_module_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
xor_module xor_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
xor_module xor_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
xor_module xor_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
xor_module xor_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
mux_module mux_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
mux_module mux_module_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
xor_module xor_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
mux_module mux_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
xor_module xor_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
xor_module xor_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
xor_module xor_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
xor_module xor_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
xor_module xor_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
xor_module xor_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
mux_module mux_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
mux_module mux_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
xor_module xor_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
xor_module xor_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
xor_module xor_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
xor_module xor_module_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
xor_module xor_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
mux_module mux_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
xor_module xor_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
xor_module xor_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
xor_module xor_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
xor_module xor_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
mux_module mux_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
xor_module xor_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
xor_module xor_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
mux_module mux_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
xor_module xor_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
mux_module mux_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
mux_module mux_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
mux_module mux_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
xor_module xor_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
xor_module xor_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
xor_module xor_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
xor_module xor_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
xor_module xor_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
xor_module xor_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
mux_module mux_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
xor_module xor_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
xor_module xor_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
xor_module xor_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
xor_module xor_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
xor_module xor_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
xor_module xor_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
xor_module xor_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
xor_module xor_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
mux_module mux_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
xor_module xor_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
xor_module xor_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
xor_module xor_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
xor_module xor_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
mux_module mux_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
xor_module xor_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
xor_module xor_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
xor_module xor_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640])); 
xor_module xor_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
xor_module xor_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
xor_module xor_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
xor_module xor_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
xor_module xor_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
mux_module mux_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
mux_module mux_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
mux_module mux_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
mux_module mux_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
xor_module xor_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
xor_module xor_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
mux_module mux_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
mux_module mux_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
xor_module xor_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
mux_module mux_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
xor_module xor_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
mux_module mux_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
xor_module xor_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
xor_module xor_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
mux_module mux_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
mux_module mux_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
xor_module xor_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
mux_module mux_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
xor_module xor_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
mux_module mux_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
mux_module mux_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
xor_module xor_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
xor_module xor_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
mux_module mux_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
xor_module xor_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
xor_module xor_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
mux_module mux_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
xor_module xor_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
mux_module mux_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
xor_module xor_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
mux_module mux_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
mux_module mux_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
mux_module mux_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
xor_module xor_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
xor_module xor_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
mux_module mux_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
xor_module xor_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
xor_module xor_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
xor_module xor_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
xor_module xor_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
xor_module xor_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
mux_module mux_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
xor_module xor_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
xor_module xor_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
xor_module xor_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
xor_module xor_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
mux_module mux_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
xor_module xor_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
mux_module mux_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
mux_module mux_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
xor_module xor_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
xor_module xor_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
mux_module mux_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
xor_module xor_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
xor_module xor_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
xor_module xor_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
xor_module xor_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
mux_module mux_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
xor_module xor_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
mux_module mux_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
xor_module xor_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
xor_module xor_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
xor_module xor_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
xor_module xor_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
xor_module xor_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
xor_module xor_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
mux_module mux_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
xor_module xor_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
mux_module mux_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
mux_module mux_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
mux_module mux_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
mux_module mux_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
mux_module mux_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
mux_module mux_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
mux_module mux_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
xor_module xor_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
xor_module xor_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
xor_module xor_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
xor_module xor_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
mux_module mux_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
xor_module xor_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
xor_module xor_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
mux_module mux_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
xor_module xor_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
xor_module xor_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
xor_module xor_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
xor_module xor_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
xor_module xor_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
xor_module xor_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
mux_module mux_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
mux_module mux_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
xor_module xor_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
xor_module xor_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
mux_module mux_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
xor_module xor_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
xor_module xor_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
xor_module xor_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
mux_module mux_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
xor_module xor_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
mux_module mux_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
xor_module xor_module_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
xor_module xor_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
xor_module xor_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
xor_module xor_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
mux_module mux_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
mux_module mux_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
xor_module xor_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
xor_module xor_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
xor_module xor_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
xor_module xor_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
xor_module xor_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
mux_module mux_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
mux_module mux_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
mux_module mux_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
xor_module xor_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
mux_module mux_module_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
mux_module mux_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
xor_module xor_module_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
xor_module xor_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
mux_module mux_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
xor_module xor_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
xor_module xor_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
xor_module xor_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
xor_module xor_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
xor_module xor_module_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
mux_module mux_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
mux_module mux_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
mux_module mux_module_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
mux_module mux_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
mux_module mux_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
mux_module mux_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
mux_module mux_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
mux_module mux_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
xor_module xor_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
mux_module mux_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
mux_module mux_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
xor_module xor_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
xor_module xor_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
mux_module mux_module_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
xor_module xor_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
mux_module mux_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
xor_module xor_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
xor_module xor_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
mux_module mux_module_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
mux_module mux_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
xor_module xor_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
mux_module mux_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
xor_module xor_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
mux_module mux_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
xor_module xor_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
mux_module mux_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
mux_module mux_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
xor_module xor_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
mux_module mux_module_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
xor_module xor_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
xor_module xor_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
mux_module mux_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
xor_module xor_module_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
mux_module mux_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
xor_module xor_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
xor_module xor_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
mux_module mux_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
xor_module xor_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
xor_module xor_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
mux_module mux_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
xor_module xor_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
xor_module xor_module_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
mux_module mux_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
mux_module mux_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
mux_module mux_module_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
xor_module xor_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
xor_module xor_module_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
xor_module xor_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
mux_module mux_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
xor_module xor_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
mux_module mux_module_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
mux_module mux_module_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
mux_module mux_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
mux_module mux_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
mux_module mux_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
xor_module xor_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
mux_module mux_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
xor_module xor_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
xor_module xor_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
xor_module xor_module_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
xor_module xor_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
xor_module xor_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
xor_module xor_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
xor_module xor_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
xor_module xor_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
mux_module mux_module_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
mux_module mux_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
mux_module mux_module_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
xor_module xor_module_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
xor_module xor_module_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
xor_module xor_module_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
mux_module mux_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
mux_module mux_module_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
xor_module xor_module_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
mux_module mux_module_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
mux_module mux_module_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
xor_module xor_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
mux_module mux_module_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
xor_module xor_module_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
xor_module xor_module_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
xor_module xor_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
xor_module xor_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
mux_module mux_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
xor_module xor_module_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
mux_module mux_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
mux_module mux_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
mux_module mux_module_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
xor_module xor_module_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
xor_module xor_module_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
mux_module mux_module_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
mux_module mux_module_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
xor_module xor_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
xor_module xor_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
mux_module mux_module_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
xor_module xor_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
xor_module xor_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
mux_module mux_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
xor_module xor_module_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
xor_module xor_module_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
xor_module xor_module_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
mux_module mux_module_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
xor_module xor_module_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
mux_module mux_module_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
xor_module xor_module_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
mux_module mux_module_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
xor_module xor_module_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
xor_module xor_module_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
xor_module xor_module_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
xor_module xor_module_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
xor_module xor_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
xor_module xor_module_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
xor_module xor_module_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
mux_module mux_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
mux_module mux_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
mux_module mux_module_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
mux_module mux_module_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
mux_module mux_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
mux_module mux_module_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
mux_module mux_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
mux_module mux_module_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
mux_module mux_module_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
xor_module xor_module_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
xor_module xor_module_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
xor_module xor_module_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
mux_module mux_module_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
xor_module xor_module_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
mux_module mux_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
mux_module mux_module_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
mux_module mux_module_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
xor_module xor_module_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
xor_module xor_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
mux_module mux_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
xor_module xor_module_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
mux_module mux_module_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
xor_module xor_module_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
mux_module mux_module_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
xor_module xor_module_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
xor_module xor_module_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
mux_module mux_module_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
xor_module xor_module_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
mux_module mux_module_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
mux_module mux_module_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
mux_module mux_module_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
xor_module xor_module_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
mux_module mux_module_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
mux_module mux_module_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
xor_module xor_module_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
mux_module mux_module_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
xor_module xor_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
xor_module xor_module_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
reg [671:0]intermediate_reg_2; 
 
mux_module mux_module_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1343]),.i2(intermediate_reg_1[1342]),.o(intermediate_reg_2[671]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1341]),.i2(intermediate_reg_1[1340]),.o(intermediate_reg_2[670]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1339]),.i2(intermediate_reg_1[1338]),.o(intermediate_reg_2[669]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1337]),.i2(intermediate_reg_1[1336]),.o(intermediate_reg_2[668]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1335]),.i2(intermediate_reg_1[1334]),.o(intermediate_reg_2[667]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1333]),.i2(intermediate_reg_1[1332]),.o(intermediate_reg_2[666]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1331]),.i2(intermediate_reg_1[1330]),.o(intermediate_reg_2[665])); 
mux_module mux_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1329]),.i2(intermediate_reg_1[1328]),.o(intermediate_reg_2[664]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1327]),.i2(intermediate_reg_1[1326]),.o(intermediate_reg_2[663])); 
mux_module mux_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1325]),.i2(intermediate_reg_1[1324]),.o(intermediate_reg_2[662]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1323]),.i2(intermediate_reg_1[1322]),.o(intermediate_reg_2[661])); 
xor_module xor_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1321]),.i2(intermediate_reg_1[1320]),.o(intermediate_reg_2[660])); 
xor_module xor_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1319]),.i2(intermediate_reg_1[1318]),.o(intermediate_reg_2[659])); 
mux_module mux_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1317]),.i2(intermediate_reg_1[1316]),.o(intermediate_reg_2[658]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1315]),.i2(intermediate_reg_1[1314]),.o(intermediate_reg_2[657]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1313]),.i2(intermediate_reg_1[1312]),.o(intermediate_reg_2[656])); 
xor_module xor_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1311]),.i2(intermediate_reg_1[1310]),.o(intermediate_reg_2[655])); 
mux_module mux_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1309]),.i2(intermediate_reg_1[1308]),.o(intermediate_reg_2[654]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1307]),.i2(intermediate_reg_1[1306]),.o(intermediate_reg_2[653])); 
mux_module mux_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1305]),.i2(intermediate_reg_1[1304]),.o(intermediate_reg_2[652]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1303]),.i2(intermediate_reg_1[1302]),.o(intermediate_reg_2[651]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1301]),.i2(intermediate_reg_1[1300]),.o(intermediate_reg_2[650]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1299]),.i2(intermediate_reg_1[1298]),.o(intermediate_reg_2[649])); 
mux_module mux_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1297]),.i2(intermediate_reg_1[1296]),.o(intermediate_reg_2[648]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1295]),.i2(intermediate_reg_1[1294]),.o(intermediate_reg_2[647]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1293]),.i2(intermediate_reg_1[1292]),.o(intermediate_reg_2[646]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1291]),.i2(intermediate_reg_1[1290]),.o(intermediate_reg_2[645])); 
mux_module mux_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1289]),.i2(intermediate_reg_1[1288]),.o(intermediate_reg_2[644]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1287]),.i2(intermediate_reg_1[1286]),.o(intermediate_reg_2[643]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1285]),.i2(intermediate_reg_1[1284]),.o(intermediate_reg_2[642]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1283]),.i2(intermediate_reg_1[1282]),.o(intermediate_reg_2[641])); 
mux_module mux_module_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1281]),.i2(intermediate_reg_1[1280]),.o(intermediate_reg_2[640]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1279]),.i2(intermediate_reg_1[1278]),.o(intermediate_reg_2[639]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1277]),.i2(intermediate_reg_1[1276]),.o(intermediate_reg_2[638]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1275]),.i2(intermediate_reg_1[1274]),.o(intermediate_reg_2[637]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1273]),.i2(intermediate_reg_1[1272]),.o(intermediate_reg_2[636]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1271]),.i2(intermediate_reg_1[1270]),.o(intermediate_reg_2[635])); 
mux_module mux_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1269]),.i2(intermediate_reg_1[1268]),.o(intermediate_reg_2[634]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1267]),.i2(intermediate_reg_1[1266]),.o(intermediate_reg_2[633]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1265]),.i2(intermediate_reg_1[1264]),.o(intermediate_reg_2[632])); 
mux_module mux_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1263]),.i2(intermediate_reg_1[1262]),.o(intermediate_reg_2[631]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1261]),.i2(intermediate_reg_1[1260]),.o(intermediate_reg_2[630])); 
xor_module xor_module_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1259]),.i2(intermediate_reg_1[1258]),.o(intermediate_reg_2[629])); 
xor_module xor_module_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1257]),.i2(intermediate_reg_1[1256]),.o(intermediate_reg_2[628])); 
xor_module xor_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1255]),.i2(intermediate_reg_1[1254]),.o(intermediate_reg_2[627])); 
xor_module xor_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1253]),.i2(intermediate_reg_1[1252]),.o(intermediate_reg_2[626])); 
xor_module xor_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1251]),.i2(intermediate_reg_1[1250]),.o(intermediate_reg_2[625])); 
xor_module xor_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1249]),.i2(intermediate_reg_1[1248]),.o(intermediate_reg_2[624])); 
mux_module mux_module_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1247]),.i2(intermediate_reg_1[1246]),.o(intermediate_reg_2[623]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1245]),.i2(intermediate_reg_1[1244]),.o(intermediate_reg_2[622]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1243]),.i2(intermediate_reg_1[1242]),.o(intermediate_reg_2[621]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1241]),.i2(intermediate_reg_1[1240]),.o(intermediate_reg_2[620])); 
xor_module xor_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1239]),.i2(intermediate_reg_1[1238]),.o(intermediate_reg_2[619])); 
mux_module mux_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1237]),.i2(intermediate_reg_1[1236]),.o(intermediate_reg_2[618]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1235]),.i2(intermediate_reg_1[1234]),.o(intermediate_reg_2[617]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1233]),.i2(intermediate_reg_1[1232]),.o(intermediate_reg_2[616])); 
mux_module mux_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1231]),.i2(intermediate_reg_1[1230]),.o(intermediate_reg_2[615]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1229]),.i2(intermediate_reg_1[1228]),.o(intermediate_reg_2[614]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1227]),.i2(intermediate_reg_1[1226]),.o(intermediate_reg_2[613]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1225]),.i2(intermediate_reg_1[1224]),.o(intermediate_reg_2[612]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1223]),.i2(intermediate_reg_1[1222]),.o(intermediate_reg_2[611])); 
mux_module mux_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1221]),.i2(intermediate_reg_1[1220]),.o(intermediate_reg_2[610]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1219]),.i2(intermediate_reg_1[1218]),.o(intermediate_reg_2[609]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1217]),.i2(intermediate_reg_1[1216]),.o(intermediate_reg_2[608])); 
xor_module xor_module_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1215]),.i2(intermediate_reg_1[1214]),.o(intermediate_reg_2[607])); 
xor_module xor_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1213]),.i2(intermediate_reg_1[1212]),.o(intermediate_reg_2[606])); 
mux_module mux_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1211]),.i2(intermediate_reg_1[1210]),.o(intermediate_reg_2[605]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1209]),.i2(intermediate_reg_1[1208]),.o(intermediate_reg_2[604])); 
xor_module xor_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1207]),.i2(intermediate_reg_1[1206]),.o(intermediate_reg_2[603])); 
mux_module mux_module_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1205]),.i2(intermediate_reg_1[1204]),.o(intermediate_reg_2[602]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1203]),.i2(intermediate_reg_1[1202]),.o(intermediate_reg_2[601]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1201]),.i2(intermediate_reg_1[1200]),.o(intermediate_reg_2[600]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1199]),.i2(intermediate_reg_1[1198]),.o(intermediate_reg_2[599])); 
mux_module mux_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1197]),.i2(intermediate_reg_1[1196]),.o(intermediate_reg_2[598]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1195]),.i2(intermediate_reg_1[1194]),.o(intermediate_reg_2[597])); 
mux_module mux_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1193]),.i2(intermediate_reg_1[1192]),.o(intermediate_reg_2[596]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1191]),.i2(intermediate_reg_1[1190]),.o(intermediate_reg_2[595])); 
mux_module mux_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1189]),.i2(intermediate_reg_1[1188]),.o(intermediate_reg_2[594]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1187]),.i2(intermediate_reg_1[1186]),.o(intermediate_reg_2[593])); 
mux_module mux_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1185]),.i2(intermediate_reg_1[1184]),.o(intermediate_reg_2[592]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1183]),.i2(intermediate_reg_1[1182]),.o(intermediate_reg_2[591])); 
mux_module mux_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1181]),.i2(intermediate_reg_1[1180]),.o(intermediate_reg_2[590]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1179]),.i2(intermediate_reg_1[1178]),.o(intermediate_reg_2[589]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1177]),.i2(intermediate_reg_1[1176]),.o(intermediate_reg_2[588])); 
mux_module mux_module_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1175]),.i2(intermediate_reg_1[1174]),.o(intermediate_reg_2[587]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1173]),.i2(intermediate_reg_1[1172]),.o(intermediate_reg_2[586])); 
xor_module xor_module_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1171]),.i2(intermediate_reg_1[1170]),.o(intermediate_reg_2[585])); 
xor_module xor_module_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1169]),.i2(intermediate_reg_1[1168]),.o(intermediate_reg_2[584])); 
xor_module xor_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1167]),.i2(intermediate_reg_1[1166]),.o(intermediate_reg_2[583])); 
xor_module xor_module_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1165]),.i2(intermediate_reg_1[1164]),.o(intermediate_reg_2[582])); 
xor_module xor_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1163]),.i2(intermediate_reg_1[1162]),.o(intermediate_reg_2[581])); 
mux_module mux_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1161]),.i2(intermediate_reg_1[1160]),.o(intermediate_reg_2[580]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1159]),.i2(intermediate_reg_1[1158]),.o(intermediate_reg_2[579]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1157]),.i2(intermediate_reg_1[1156]),.o(intermediate_reg_2[578])); 
xor_module xor_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1155]),.i2(intermediate_reg_1[1154]),.o(intermediate_reg_2[577])); 
mux_module mux_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1153]),.i2(intermediate_reg_1[1152]),.o(intermediate_reg_2[576]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1151]),.i2(intermediate_reg_1[1150]),.o(intermediate_reg_2[575]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1149]),.i2(intermediate_reg_1[1148]),.o(intermediate_reg_2[574]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1147]),.i2(intermediate_reg_1[1146]),.o(intermediate_reg_2[573])); 
mux_module mux_module_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1145]),.i2(intermediate_reg_1[1144]),.o(intermediate_reg_2[572]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1143]),.i2(intermediate_reg_1[1142]),.o(intermediate_reg_2[571])); 
xor_module xor_module_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1141]),.i2(intermediate_reg_1[1140]),.o(intermediate_reg_2[570])); 
xor_module xor_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1139]),.i2(intermediate_reg_1[1138]),.o(intermediate_reg_2[569])); 
mux_module mux_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1137]),.i2(intermediate_reg_1[1136]),.o(intermediate_reg_2[568]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1135]),.i2(intermediate_reg_1[1134]),.o(intermediate_reg_2[567]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1133]),.i2(intermediate_reg_1[1132]),.o(intermediate_reg_2[566])); 
xor_module xor_module_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1131]),.i2(intermediate_reg_1[1130]),.o(intermediate_reg_2[565])); 
xor_module xor_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1129]),.i2(intermediate_reg_1[1128]),.o(intermediate_reg_2[564])); 
mux_module mux_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1127]),.i2(intermediate_reg_1[1126]),.o(intermediate_reg_2[563]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1125]),.i2(intermediate_reg_1[1124]),.o(intermediate_reg_2[562])); 
xor_module xor_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1123]),.i2(intermediate_reg_1[1122]),.o(intermediate_reg_2[561])); 
mux_module mux_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1121]),.i2(intermediate_reg_1[1120]),.o(intermediate_reg_2[560]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1119]),.i2(intermediate_reg_1[1118]),.o(intermediate_reg_2[559]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1117]),.i2(intermediate_reg_1[1116]),.o(intermediate_reg_2[558])); 
xor_module xor_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1115]),.i2(intermediate_reg_1[1114]),.o(intermediate_reg_2[557])); 
mux_module mux_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1113]),.i2(intermediate_reg_1[1112]),.o(intermediate_reg_2[556]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1111]),.i2(intermediate_reg_1[1110]),.o(intermediate_reg_2[555]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1109]),.i2(intermediate_reg_1[1108]),.o(intermediate_reg_2[554]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1107]),.i2(intermediate_reg_1[1106]),.o(intermediate_reg_2[553]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1105]),.i2(intermediate_reg_1[1104]),.o(intermediate_reg_2[552])); 
xor_module xor_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1103]),.i2(intermediate_reg_1[1102]),.o(intermediate_reg_2[551])); 
xor_module xor_module_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1101]),.i2(intermediate_reg_1[1100]),.o(intermediate_reg_2[550])); 
xor_module xor_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1099]),.i2(intermediate_reg_1[1098]),.o(intermediate_reg_2[549])); 
mux_module mux_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1097]),.i2(intermediate_reg_1[1096]),.o(intermediate_reg_2[548]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1095]),.i2(intermediate_reg_1[1094]),.o(intermediate_reg_2[547]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1093]),.i2(intermediate_reg_1[1092]),.o(intermediate_reg_2[546]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1091]),.i2(intermediate_reg_1[1090]),.o(intermediate_reg_2[545])); 
mux_module mux_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1089]),.i2(intermediate_reg_1[1088]),.o(intermediate_reg_2[544]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1087]),.i2(intermediate_reg_1[1086]),.o(intermediate_reg_2[543])); 
mux_module mux_module_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1085]),.i2(intermediate_reg_1[1084]),.o(intermediate_reg_2[542]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1083]),.i2(intermediate_reg_1[1082]),.o(intermediate_reg_2[541]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1081]),.i2(intermediate_reg_1[1080]),.o(intermediate_reg_2[540])); 
xor_module xor_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1079]),.i2(intermediate_reg_1[1078]),.o(intermediate_reg_2[539])); 
xor_module xor_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1077]),.i2(intermediate_reg_1[1076]),.o(intermediate_reg_2[538])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1075]),.i2(intermediate_reg_1[1074]),.o(intermediate_reg_2[537]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1073]),.i2(intermediate_reg_1[1072]),.o(intermediate_reg_2[536]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1071]),.i2(intermediate_reg_1[1070]),.o(intermediate_reg_2[535])); 
mux_module mux_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1069]),.i2(intermediate_reg_1[1068]),.o(intermediate_reg_2[534]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1067]),.i2(intermediate_reg_1[1066]),.o(intermediate_reg_2[533])); 
mux_module mux_module_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1065]),.i2(intermediate_reg_1[1064]),.o(intermediate_reg_2[532]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1063]),.i2(intermediate_reg_1[1062]),.o(intermediate_reg_2[531])); 
xor_module xor_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1061]),.i2(intermediate_reg_1[1060]),.o(intermediate_reg_2[530])); 
xor_module xor_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1059]),.i2(intermediate_reg_1[1058]),.o(intermediate_reg_2[529])); 
mux_module mux_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1057]),.i2(intermediate_reg_1[1056]),.o(intermediate_reg_2[528]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1055]),.i2(intermediate_reg_1[1054]),.o(intermediate_reg_2[527])); 
mux_module mux_module_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1053]),.i2(intermediate_reg_1[1052]),.o(intermediate_reg_2[526]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1051]),.i2(intermediate_reg_1[1050]),.o(intermediate_reg_2[525]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1049]),.i2(intermediate_reg_1[1048]),.o(intermediate_reg_2[524])); 
mux_module mux_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1047]),.i2(intermediate_reg_1[1046]),.o(intermediate_reg_2[523]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1045]),.i2(intermediate_reg_1[1044]),.o(intermediate_reg_2[522])); 
xor_module xor_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1043]),.i2(intermediate_reg_1[1042]),.o(intermediate_reg_2[521])); 
mux_module mux_module_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1041]),.i2(intermediate_reg_1[1040]),.o(intermediate_reg_2[520]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1039]),.i2(intermediate_reg_1[1038]),.o(intermediate_reg_2[519])); 
mux_module mux_module_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1037]),.i2(intermediate_reg_1[1036]),.o(intermediate_reg_2[518]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1035]),.i2(intermediate_reg_1[1034]),.o(intermediate_reg_2[517])); 
mux_module mux_module_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1033]),.i2(intermediate_reg_1[1032]),.o(intermediate_reg_2[516]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1031]),.i2(intermediate_reg_1[1030]),.o(intermediate_reg_2[515]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1029]),.i2(intermediate_reg_1[1028]),.o(intermediate_reg_2[514])); 
xor_module xor_module_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513])); 
xor_module xor_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512])); 
xor_module xor_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511])); 
xor_module xor_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510])); 
mux_module mux_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508])); 
xor_module xor_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507])); 
xor_module xor_module_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506])); 
mux_module mux_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504])); 
xor_module xor_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503])); 
mux_module mux_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499])); 
xor_module xor_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498])); 
mux_module mux_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495])); 
xor_module xor_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494])); 
mux_module mux_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491])); 
xor_module xor_module_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490])); 
xor_module xor_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489])); 
mux_module mux_module_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487])); 
mux_module mux_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485])); 
mux_module mux_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482])); 
mux_module mux_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
mux_module mux_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475])); 
xor_module xor_module_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474])); 
mux_module mux_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472])); 
xor_module xor_module_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471])); 
mux_module mux_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469])); 
mux_module mux_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467])); 
mux_module mux_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465])); 
mux_module mux_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463])); 
xor_module xor_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462])); 
mux_module mux_module_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460])); 
mux_module mux_module_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457])); 
xor_module xor_module_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456])); 
xor_module xor_module_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455])); 
mux_module mux_module_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453])); 
mux_module mux_module_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450])); 
xor_module xor_module_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449])); 
mux_module mux_module_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445])); 
mux_module mux_module_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443])); 
xor_module xor_module_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442])); 
mux_module mux_module_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435])); 
xor_module xor_module_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434])); 
mux_module mux_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429])); 
xor_module xor_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428])); 
xor_module xor_module_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427])); 
xor_module xor_module_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426])); 
mux_module mux_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424])); 
mux_module mux_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420])); 
xor_module xor_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419])); 
mux_module mux_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417])); 
xor_module xor_module_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416])); 
mux_module mux_module_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414])); 
xor_module xor_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413])); 
xor_module xor_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412])); 
xor_module xor_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411])); 
xor_module xor_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410])); 
mux_module mux_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407])); 
mux_module mux_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404])); 
xor_module xor_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403])); 
mux_module mux_module_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401])); 
xor_module xor_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400])); 
xor_module xor_module_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399])); 
mux_module mux_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397])); 
xor_module xor_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396])); 
xor_module xor_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395])); 
mux_module mux_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393])); 
mux_module mux_module_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389])); 
xor_module xor_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388])); 
mux_module mux_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386])); 
mux_module mux_module_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384])); 
mux_module mux_module_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
xor_module xor_module_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
xor_module xor_module_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379])); 
mux_module mux_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375])); 
mux_module mux_module_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372])); 
mux_module mux_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
mux_module mux_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368])); 
mux_module mux_module_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366])); 
xor_module xor_module_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365])); 
xor_module xor_module_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
mux_module mux_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362])); 
mux_module mux_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360])); 
xor_module xor_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
mux_module mux_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354])); 
mux_module mux_module_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352])); 
xor_module xor_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351])); 
mux_module mux_module_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348])); 
xor_module xor_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
mux_module mux_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
mux_module mux_module_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342])); 
xor_module xor_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341])); 
xor_module xor_module_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340])); 
xor_module xor_module_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339])); 
mux_module mux_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336])); 
xor_module xor_module_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
xor_module xor_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334])); 
xor_module xor_module_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333])); 
xor_module xor_module_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332])); 
mux_module mux_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
xor_module xor_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
xor_module xor_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328])); 
xor_module xor_module_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
xor_module xor_module_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326])); 
xor_module xor_module_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325])); 
mux_module mux_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318])); 
mux_module mux_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315])); 
xor_module xor_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314])); 
mux_module mux_module_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312])); 
xor_module xor_module_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311])); 
mux_module mux_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307])); 
xor_module xor_module_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306])); 
mux_module mux_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302])); 
xor_module xor_module_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
mux_module mux_module_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299])); 
xor_module xor_module_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298])); 
mux_module mux_module_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
mux_module mux_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292])); 
xor_module xor_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291])); 
mux_module mux_module_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288])); 
mux_module mux_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
mux_module mux_module_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
mux_module mux_module_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280])); 
mux_module mux_module_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
xor_module xor_module_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
xor_module xor_module_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
xor_module xor_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
xor_module xor_module_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270])); 
xor_module xor_module_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
mux_module mux_module_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
xor_module xor_module_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264])); 
xor_module xor_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263])); 
xor_module xor_module_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
xor_module xor_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261])); 
mux_module mux_module_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258])); 
xor_module xor_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257])); 
mux_module mux_module_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
xor_module xor_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250])); 
xor_module xor_module_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
mux_module mux_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246])); 
xor_module xor_module_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
mux_module mux_module_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
xor_module xor_module_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240])); 
mux_module mux_module_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
mux_module mux_module_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235])); 
xor_module xor_module_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
mux_module mux_module_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229])); 
xor_module xor_module_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
mux_module mux_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
mux_module mux_module_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223])); 
xor_module xor_module_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
mux_module mux_module_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220])); 
mux_module mux_module_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215])); 
mux_module mux_module_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
mux_module mux_module_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209])); 
mux_module mux_module_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
xor_module xor_module_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
xor_module xor_module_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
xor_module xor_module_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204])); 
mux_module mux_module_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202])); 
xor_module xor_module_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201])); 
mux_module mux_module_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
xor_module xor_module_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198])); 
mux_module mux_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193])); 
xor_module xor_module_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
xor_module xor_module_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
mux_module mux_module_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186])); 
mux_module mux_module_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
xor_module xor_module_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183])); 
mux_module mux_module_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180])); 
mux_module mux_module_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178])); 
mux_module mux_module_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
mux_module mux_module_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
xor_module xor_module_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
mux_module mux_module_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
xor_module xor_module_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164])); 
xor_module xor_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
mux_module mux_module_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160])); 
xor_module xor_module_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
xor_module xor_module_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158])); 
mux_module mux_module_inst_2_514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154])); 
xor_module xor_module_inst_2_518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153])); 
mux_module mux_module_inst_2_519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
mux_module mux_module_inst_2_523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146])); 
xor_module xor_module_inst_2_526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145])); 
xor_module xor_module_inst_2_527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144])); 
mux_module mux_module_inst_2_528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140])); 
mux_module mux_module_inst_2_532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
xor_module xor_module_inst_2_535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136])); 
xor_module xor_module_inst_2_536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135])); 
mux_module mux_module_inst_2_537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129])); 
mux_module mux_module_inst_2_543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
xor_module xor_module_inst_2_547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124])); 
mux_module mux_module_inst_2_548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
mux_module mux_module_inst_2_550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119])); 
mux_module mux_module_inst_2_553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113])); 
mux_module mux_module_inst_2_559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_560(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111])); 
xor_module xor_module_inst_2_561(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
xor_module xor_module_inst_2_562(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
xor_module xor_module_inst_2_563(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
xor_module xor_module_inst_2_564(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107])); 
xor_module xor_module_inst_2_565(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
mux_module mux_module_inst_2_566(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_567(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104])); 
xor_module xor_module_inst_2_568(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
mux_module mux_module_inst_2_569(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_570(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
xor_module xor_module_inst_2_571(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100])); 
mux_module mux_module_inst_2_572(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_573(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98])); 
xor_module xor_module_inst_2_574(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
mux_module mux_module_inst_2_575(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_576(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_577(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_578(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
mux_module mux_module_inst_2_579(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_580(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_581(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_582(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89])); 
xor_module xor_module_inst_2_583(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88])); 
xor_module xor_module_inst_2_584(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
mux_module mux_module_inst_2_585(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_586(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
xor_module xor_module_inst_2_587(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
mux_module mux_module_inst_2_588(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_589(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_590(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
xor_module xor_module_inst_2_591(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80])); 
xor_module xor_module_inst_2_592(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79])); 
mux_module mux_module_inst_2_593(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_594(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
mux_module mux_module_inst_2_595(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_596(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_597(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74])); 
mux_module mux_module_inst_2_598(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_599(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72])); 
mux_module mux_module_inst_2_600(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_601(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
mux_module mux_module_inst_2_602(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_603(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_604(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_605(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_606(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65])); 
xor_module xor_module_inst_2_607(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64])); 
xor_module xor_module_inst_2_608(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
xor_module xor_module_inst_2_609(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
xor_module xor_module_inst_2_610(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
mux_module mux_module_inst_2_611(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_612(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_613(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_614(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_615(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56])); 
mux_module mux_module_inst_2_616(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_617(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_618(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
xor_module xor_module_inst_2_619(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
xor_module xor_module_inst_2_620(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51])); 
xor_module xor_module_inst_2_621(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
xor_module xor_module_inst_2_622(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
mux_module mux_module_inst_2_623(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_624(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_625(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_626(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_627(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_628(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
mux_module mux_module_inst_2_629(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_630(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_631(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_632(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_633(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_634(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
xor_module xor_module_inst_2_635(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36])); 
xor_module xor_module_inst_2_636(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35])); 
mux_module mux_module_inst_2_637(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_638(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_639(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_640(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_641(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_642(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_643(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_644(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_645(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_646(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25])); 
xor_module xor_module_inst_2_647(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
xor_module xor_module_inst_2_648(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23])); 
mux_module mux_module_inst_2_649(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_650(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_651(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_652(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
xor_module xor_module_inst_2_653(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18])); 
mux_module mux_module_inst_2_654(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_655(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
xor_module xor_module_inst_2_656(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15])); 
mux_module mux_module_inst_2_657(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_658(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_659(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_660(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_661(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_662(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
mux_module mux_module_inst_2_663(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_664(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
mux_module mux_module_inst_2_665(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_666(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5])); 
xor_module xor_module_inst_2_667(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
xor_module xor_module_inst_2_668(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
mux_module mux_module_inst_2_669(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_670(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
mux_module mux_module_inst_2_671(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0]),.sel(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [671:0] <= intermediate_reg_2; 
outp[1055:672] <= intermediate_reg_2[383:0] ; 
end 
endmodule 
 

module interface_15(input [975:0] inp, output reg [1253:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[975:0] <= inp ; 
outp[1253:976] <= inp[277:0] ; 
end 
endmodule 

module interface_16(input [127:0] inp, output reg [417:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[127:0] <= inp ; 
outp[255:128] <= inp ; 
outp[383:256] <= inp ; 
outp[417:384] <= inp[33:0] ; 
end 
endmodule 

module interface_17(input [287:0] inp, output reg [1271:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[287:0] <= inp ; 
outp[575:288] <= inp ; 
outp[863:576] <= inp ; 
outp[1151:864] <= inp ; 
outp[1271:1152] <= inp[119:0] ; 
end 
endmodule 

module interface_18(input [959:0] inp, output reg [794:0] outp, input clk, input reset);
reg [959:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [479:0]intermediate_reg_1; 
 
xor_module xor_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
xor_module xor_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
xor_module xor_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
xor_module xor_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
xor_module xor_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
xor_module xor_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
xor_module xor_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
xor_module xor_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
xor_module xor_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
xor_module xor_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
xor_module xor_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
mux_module mux_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
mux_module mux_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
xor_module xor_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
xor_module xor_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
xor_module xor_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
xor_module xor_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
xor_module xor_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
xor_module xor_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
xor_module xor_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
xor_module xor_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
xor_module xor_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
xor_module xor_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
xor_module xor_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
xor_module xor_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
mux_module mux_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
xor_module xor_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
mux_module mux_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
xor_module xor_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
xor_module xor_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
xor_module xor_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
xor_module xor_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
xor_module xor_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
xor_module xor_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
xor_module xor_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
xor_module xor_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
xor_module xor_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
mux_module mux_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
xor_module xor_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
mux_module mux_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
mux_module mux_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
xor_module xor_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
xor_module xor_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
mux_module mux_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
xor_module xor_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
xor_module xor_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
xor_module xor_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
xor_module xor_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
xor_module xor_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
xor_module xor_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
xor_module xor_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
xor_module xor_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
xor_module xor_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
xor_module xor_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
xor_module xor_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
xor_module xor_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
xor_module xor_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
mux_module mux_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
xor_module xor_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
mux_module mux_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
xor_module xor_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
xor_module xor_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
xor_module xor_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
xor_module xor_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
xor_module xor_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
xor_module xor_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
xor_module xor_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
xor_module xor_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
xor_module xor_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
mux_module mux_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
mux_module mux_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
xor_module xor_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
xor_module xor_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
xor_module xor_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
mux_module mux_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
mux_module mux_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
xor_module xor_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
mux_module mux_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
mux_module mux_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
xor_module xor_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
xor_module xor_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
xor_module xor_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
mux_module mux_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
xor_module xor_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
xor_module xor_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
xor_module xor_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
xor_module xor_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
xor_module xor_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
xor_module xor_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
mux_module mux_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
xor_module xor_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
xor_module xor_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
xor_module xor_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
xor_module xor_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
xor_module xor_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
mux_module mux_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
xor_module xor_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
xor_module xor_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
xor_module xor_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
xor_module xor_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
xor_module xor_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
xor_module xor_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
xor_module xor_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
mux_module mux_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
xor_module xor_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
mux_module mux_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
xor_module xor_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
xor_module xor_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
mux_module mux_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
xor_module xor_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
mux_module mux_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
xor_module xor_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
xor_module xor_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
xor_module xor_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
xor_module xor_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
xor_module xor_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
mux_module mux_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
xor_module xor_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
xor_module xor_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
xor_module xor_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
xor_module xor_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
xor_module xor_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
xor_module xor_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
xor_module xor_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
xor_module xor_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
xor_module xor_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
xor_module xor_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
xor_module xor_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
always@(posedge clk) begin 
outp [479:0] <= intermediate_reg_1; 
outp[794:480] <= intermediate_reg_1[314:0] ; 
end 
endmodule 
 

module interface_19(input [815:0] inp, output reg [103:0] outp, input clk, input reset);
reg [815:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [407:0]intermediate_reg_1; 
 
xor_module xor_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
mux_module mux_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
mux_module mux_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
xor_module xor_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
xor_module xor_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
xor_module xor_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
xor_module xor_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
xor_module xor_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
xor_module xor_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
xor_module xor_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
xor_module xor_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
xor_module xor_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
xor_module xor_module_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
xor_module xor_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
xor_module xor_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
xor_module xor_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
mux_module mux_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
xor_module xor_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
xor_module xor_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
xor_module xor_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
xor_module xor_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
xor_module xor_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
xor_module xor_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
xor_module xor_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
xor_module xor_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
mux_module mux_module_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
xor_module xor_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
mux_module mux_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
xor_module xor_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
xor_module xor_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
xor_module xor_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
xor_module xor_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
mux_module mux_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
xor_module xor_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
xor_module xor_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
xor_module xor_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
xor_module xor_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
mux_module mux_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
mux_module mux_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
xor_module xor_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
mux_module mux_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
xor_module xor_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
xor_module xor_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
xor_module xor_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
xor_module xor_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
mux_module mux_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
xor_module xor_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
xor_module xor_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
mux_module mux_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
mux_module mux_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
xor_module xor_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
xor_module xor_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
xor_module xor_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
xor_module xor_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
xor_module xor_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
xor_module xor_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
xor_module xor_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
xor_module xor_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
mux_module mux_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
xor_module xor_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
xor_module xor_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
xor_module xor_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
mux_module mux_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
xor_module xor_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
xor_module xor_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
xor_module xor_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
xor_module xor_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
mux_module mux_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
mux_module mux_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
xor_module xor_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
mux_module mux_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
xor_module xor_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
xor_module xor_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
xor_module xor_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117])); 
xor_module xor_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
xor_module xor_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115])); 
mux_module mux_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
xor_module xor_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
mux_module mux_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
xor_module xor_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
xor_module xor_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
mux_module mux_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
mux_module mux_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
xor_module xor_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
xor_module xor_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
xor_module xor_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
xor_module xor_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
mux_module mux_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
xor_module xor_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
xor_module xor_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
xor_module xor_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
xor_module xor_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
mux_module mux_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
xor_module xor_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
xor_module xor_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
xor_module xor_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
xor_module xor_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
xor_module xor_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
xor_module xor_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
xor_module xor_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
mux_module mux_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
xor_module xor_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
xor_module xor_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
xor_module xor_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
xor_module xor_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
xor_module xor_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
mux_module mux_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
mux_module mux_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
xor_module xor_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
xor_module xor_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
mux_module mux_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
xor_module xor_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
mux_module mux_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
mux_module mux_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
xor_module xor_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
xor_module xor_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
xor_module xor_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
xor_module xor_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
xor_module xor_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
xor_module xor_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
xor_module xor_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
xor_module xor_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
mux_module mux_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2]),.sel(intermediate_reg_0[0])); 
xor_module xor_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
xor_module xor_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
reg [203:0]intermediate_reg_2; 
 
xor_module xor_module_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203])); 
mux_module mux_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201])); 
mux_module mux_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
mux_module mux_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
xor_module xor_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
mux_module mux_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189])); 
xor_module xor_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
mux_module mux_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
mux_module mux_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182])); 
xor_module xor_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181])); 
mux_module mux_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
mux_module mux_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175])); 
mux_module mux_module_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
xor_module xor_module_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
mux_module mux_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
mux_module mux_module_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168])); 
mux_module mux_module_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164])); 
mux_module mux_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162])); 
mux_module mux_module_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
mux_module mux_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157])); 
mux_module mux_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154])); 
mux_module mux_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152])); 
xor_module xor_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151])); 
xor_module xor_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
xor_module xor_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
xor_module xor_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148])); 
mux_module mux_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146])); 
mux_module mux_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141])); 
xor_module xor_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140])); 
mux_module mux_module_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138])); 
xor_module xor_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
mux_module mux_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
mux_module mux_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132])); 
mux_module mux_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
xor_module xor_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
xor_module xor_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126])); 
mux_module mux_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123])); 
mux_module mux_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121])); 
mux_module mux_module_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119])); 
mux_module mux_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117])); 
mux_module mux_module_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115])); 
xor_module xor_module_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
mux_module mux_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
mux_module mux_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
xor_module xor_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
mux_module mux_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
xor_module xor_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105])); 
mux_module mux_module_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
mux_module mux_module_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
mux_module mux_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
xor_module xor_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96])); 
mux_module mux_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
mux_module mux_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
xor_module xor_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89])); 
xor_module xor_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88])); 
xor_module xor_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
xor_module xor_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
mux_module mux_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82])); 
xor_module xor_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
xor_module xor_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80])); 
mux_module mux_module_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76])); 
mux_module mux_module_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73])); 
xor_module xor_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72])); 
mux_module mux_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63])); 
xor_module xor_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
xor_module xor_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
mux_module mux_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59])); 
xor_module xor_module_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
mux_module mux_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55])); 
mux_module mux_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
mux_module mux_module_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51])); 
mux_module mux_module_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
mux_module mux_module_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
mux_module mux_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38])); 
xor_module xor_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
xor_module xor_module_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36])); 
mux_module mux_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33])); 
xor_module xor_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32])); 
xor_module xor_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
xor_module xor_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
mux_module mux_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27])); 
xor_module xor_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26])); 
xor_module xor_module_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25])); 
xor_module xor_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
mux_module mux_module_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21])); 
mux_module mux_module_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
xor_module xor_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18])); 
mux_module mux_module_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
mux_module mux_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14])); 
mux_module mux_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
xor_module xor_module_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6])); 
mux_module mux_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
xor_module xor_module_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
mux_module mux_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2]),.sel(intermediate_reg_1[0])); 
xor_module xor_module_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
mux_module mux_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0]),.sel(intermediate_reg_1[0])); 
reg [101:0]intermediate_reg_3; 
 
xor_module xor_module_inst_3_0(.clk(clk),.reset(reset),.i1(intermediate_reg_2[203]),.i2(intermediate_reg_2[202]),.o(intermediate_reg_3[101])); 
mux_module mux_module_inst_3_1(.clk(clk),.reset(reset),.i1(intermediate_reg_2[201]),.i2(intermediate_reg_2[200]),.o(intermediate_reg_3[100]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_2(.clk(clk),.reset(reset),.i1(intermediate_reg_2[199]),.i2(intermediate_reg_2[198]),.o(intermediate_reg_3[99])); 
mux_module mux_module_inst_3_3(.clk(clk),.reset(reset),.i1(intermediate_reg_2[197]),.i2(intermediate_reg_2[196]),.o(intermediate_reg_3[98]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_4(.clk(clk),.reset(reset),.i1(intermediate_reg_2[195]),.i2(intermediate_reg_2[194]),.o(intermediate_reg_3[97]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_5(.clk(clk),.reset(reset),.i1(intermediate_reg_2[193]),.i2(intermediate_reg_2[192]),.o(intermediate_reg_3[96]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_6(.clk(clk),.reset(reset),.i1(intermediate_reg_2[191]),.i2(intermediate_reg_2[190]),.o(intermediate_reg_3[95]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_7(.clk(clk),.reset(reset),.i1(intermediate_reg_2[189]),.i2(intermediate_reg_2[188]),.o(intermediate_reg_3[94])); 
xor_module xor_module_inst_3_8(.clk(clk),.reset(reset),.i1(intermediate_reg_2[187]),.i2(intermediate_reg_2[186]),.o(intermediate_reg_3[93])); 
mux_module mux_module_inst_3_9(.clk(clk),.reset(reset),.i1(intermediate_reg_2[185]),.i2(intermediate_reg_2[184]),.o(intermediate_reg_3[92]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_10(.clk(clk),.reset(reset),.i1(intermediate_reg_2[183]),.i2(intermediate_reg_2[182]),.o(intermediate_reg_3[91])); 
mux_module mux_module_inst_3_11(.clk(clk),.reset(reset),.i1(intermediate_reg_2[181]),.i2(intermediate_reg_2[180]),.o(intermediate_reg_3[90]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_12(.clk(clk),.reset(reset),.i1(intermediate_reg_2[179]),.i2(intermediate_reg_2[178]),.o(intermediate_reg_3[89])); 
mux_module mux_module_inst_3_13(.clk(clk),.reset(reset),.i1(intermediate_reg_2[177]),.i2(intermediate_reg_2[176]),.o(intermediate_reg_3[88]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_14(.clk(clk),.reset(reset),.i1(intermediate_reg_2[175]),.i2(intermediate_reg_2[174]),.o(intermediate_reg_3[87]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_15(.clk(clk),.reset(reset),.i1(intermediate_reg_2[173]),.i2(intermediate_reg_2[172]),.o(intermediate_reg_3[86])); 
mux_module mux_module_inst_3_16(.clk(clk),.reset(reset),.i1(intermediate_reg_2[171]),.i2(intermediate_reg_2[170]),.o(intermediate_reg_3[85]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_17(.clk(clk),.reset(reset),.i1(intermediate_reg_2[169]),.i2(intermediate_reg_2[168]),.o(intermediate_reg_3[84])); 
mux_module mux_module_inst_3_18(.clk(clk),.reset(reset),.i1(intermediate_reg_2[167]),.i2(intermediate_reg_2[166]),.o(intermediate_reg_3[83]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_19(.clk(clk),.reset(reset),.i1(intermediate_reg_2[165]),.i2(intermediate_reg_2[164]),.o(intermediate_reg_3[82])); 
mux_module mux_module_inst_3_20(.clk(clk),.reset(reset),.i1(intermediate_reg_2[163]),.i2(intermediate_reg_2[162]),.o(intermediate_reg_3[81]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_21(.clk(clk),.reset(reset),.i1(intermediate_reg_2[161]),.i2(intermediate_reg_2[160]),.o(intermediate_reg_3[80])); 
mux_module mux_module_inst_3_22(.clk(clk),.reset(reset),.i1(intermediate_reg_2[159]),.i2(intermediate_reg_2[158]),.o(intermediate_reg_3[79]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_23(.clk(clk),.reset(reset),.i1(intermediate_reg_2[157]),.i2(intermediate_reg_2[156]),.o(intermediate_reg_3[78]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_24(.clk(clk),.reset(reset),.i1(intermediate_reg_2[155]),.i2(intermediate_reg_2[154]),.o(intermediate_reg_3[77])); 
xor_module xor_module_inst_3_25(.clk(clk),.reset(reset),.i1(intermediate_reg_2[153]),.i2(intermediate_reg_2[152]),.o(intermediate_reg_3[76])); 
xor_module xor_module_inst_3_26(.clk(clk),.reset(reset),.i1(intermediate_reg_2[151]),.i2(intermediate_reg_2[150]),.o(intermediate_reg_3[75])); 
xor_module xor_module_inst_3_27(.clk(clk),.reset(reset),.i1(intermediate_reg_2[149]),.i2(intermediate_reg_2[148]),.o(intermediate_reg_3[74])); 
xor_module xor_module_inst_3_28(.clk(clk),.reset(reset),.i1(intermediate_reg_2[147]),.i2(intermediate_reg_2[146]),.o(intermediate_reg_3[73])); 
xor_module xor_module_inst_3_29(.clk(clk),.reset(reset),.i1(intermediate_reg_2[145]),.i2(intermediate_reg_2[144]),.o(intermediate_reg_3[72])); 
mux_module mux_module_inst_3_30(.clk(clk),.reset(reset),.i1(intermediate_reg_2[143]),.i2(intermediate_reg_2[142]),.o(intermediate_reg_3[71]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_31(.clk(clk),.reset(reset),.i1(intermediate_reg_2[141]),.i2(intermediate_reg_2[140]),.o(intermediate_reg_3[70]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_32(.clk(clk),.reset(reset),.i1(intermediate_reg_2[139]),.i2(intermediate_reg_2[138]),.o(intermediate_reg_3[69]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_33(.clk(clk),.reset(reset),.i1(intermediate_reg_2[137]),.i2(intermediate_reg_2[136]),.o(intermediate_reg_3[68]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_34(.clk(clk),.reset(reset),.i1(intermediate_reg_2[135]),.i2(intermediate_reg_2[134]),.o(intermediate_reg_3[67])); 
mux_module mux_module_inst_3_35(.clk(clk),.reset(reset),.i1(intermediate_reg_2[133]),.i2(intermediate_reg_2[132]),.o(intermediate_reg_3[66]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_36(.clk(clk),.reset(reset),.i1(intermediate_reg_2[131]),.i2(intermediate_reg_2[130]),.o(intermediate_reg_3[65])); 
mux_module mux_module_inst_3_37(.clk(clk),.reset(reset),.i1(intermediate_reg_2[129]),.i2(intermediate_reg_2[128]),.o(intermediate_reg_3[64]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_38(.clk(clk),.reset(reset),.i1(intermediate_reg_2[127]),.i2(intermediate_reg_2[126]),.o(intermediate_reg_3[63])); 
mux_module mux_module_inst_3_39(.clk(clk),.reset(reset),.i1(intermediate_reg_2[125]),.i2(intermediate_reg_2[124]),.o(intermediate_reg_3[62]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_40(.clk(clk),.reset(reset),.i1(intermediate_reg_2[123]),.i2(intermediate_reg_2[122]),.o(intermediate_reg_3[61])); 
mux_module mux_module_inst_3_41(.clk(clk),.reset(reset),.i1(intermediate_reg_2[121]),.i2(intermediate_reg_2[120]),.o(intermediate_reg_3[60]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_42(.clk(clk),.reset(reset),.i1(intermediate_reg_2[119]),.i2(intermediate_reg_2[118]),.o(intermediate_reg_3[59])); 
mux_module mux_module_inst_3_43(.clk(clk),.reset(reset),.i1(intermediate_reg_2[117]),.i2(intermediate_reg_2[116]),.o(intermediate_reg_3[58]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_44(.clk(clk),.reset(reset),.i1(intermediate_reg_2[115]),.i2(intermediate_reg_2[114]),.o(intermediate_reg_3[57]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_45(.clk(clk),.reset(reset),.i1(intermediate_reg_2[113]),.i2(intermediate_reg_2[112]),.o(intermediate_reg_3[56])); 
mux_module mux_module_inst_3_46(.clk(clk),.reset(reset),.i1(intermediate_reg_2[111]),.i2(intermediate_reg_2[110]),.o(intermediate_reg_3[55]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_47(.clk(clk),.reset(reset),.i1(intermediate_reg_2[109]),.i2(intermediate_reg_2[108]),.o(intermediate_reg_3[54])); 
mux_module mux_module_inst_3_48(.clk(clk),.reset(reset),.i1(intermediate_reg_2[107]),.i2(intermediate_reg_2[106]),.o(intermediate_reg_3[53]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_49(.clk(clk),.reset(reset),.i1(intermediate_reg_2[105]),.i2(intermediate_reg_2[104]),.o(intermediate_reg_3[52])); 
mux_module mux_module_inst_3_50(.clk(clk),.reset(reset),.i1(intermediate_reg_2[103]),.i2(intermediate_reg_2[102]),.o(intermediate_reg_3[51]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_51(.clk(clk),.reset(reset),.i1(intermediate_reg_2[101]),.i2(intermediate_reg_2[100]),.o(intermediate_reg_3[50])); 
mux_module mux_module_inst_3_52(.clk(clk),.reset(reset),.i1(intermediate_reg_2[99]),.i2(intermediate_reg_2[98]),.o(intermediate_reg_3[49]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_53(.clk(clk),.reset(reset),.i1(intermediate_reg_2[97]),.i2(intermediate_reg_2[96]),.o(intermediate_reg_3[48])); 
xor_module xor_module_inst_3_54(.clk(clk),.reset(reset),.i1(intermediate_reg_2[95]),.i2(intermediate_reg_2[94]),.o(intermediate_reg_3[47])); 
mux_module mux_module_inst_3_55(.clk(clk),.reset(reset),.i1(intermediate_reg_2[93]),.i2(intermediate_reg_2[92]),.o(intermediate_reg_3[46]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_56(.clk(clk),.reset(reset),.i1(intermediate_reg_2[91]),.i2(intermediate_reg_2[90]),.o(intermediate_reg_3[45]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_57(.clk(clk),.reset(reset),.i1(intermediate_reg_2[89]),.i2(intermediate_reg_2[88]),.o(intermediate_reg_3[44]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_58(.clk(clk),.reset(reset),.i1(intermediate_reg_2[87]),.i2(intermediate_reg_2[86]),.o(intermediate_reg_3[43])); 
xor_module xor_module_inst_3_59(.clk(clk),.reset(reset),.i1(intermediate_reg_2[85]),.i2(intermediate_reg_2[84]),.o(intermediate_reg_3[42])); 
xor_module xor_module_inst_3_60(.clk(clk),.reset(reset),.i1(intermediate_reg_2[83]),.i2(intermediate_reg_2[82]),.o(intermediate_reg_3[41])); 
mux_module mux_module_inst_3_61(.clk(clk),.reset(reset),.i1(intermediate_reg_2[81]),.i2(intermediate_reg_2[80]),.o(intermediate_reg_3[40]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_62(.clk(clk),.reset(reset),.i1(intermediate_reg_2[79]),.i2(intermediate_reg_2[78]),.o(intermediate_reg_3[39]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_63(.clk(clk),.reset(reset),.i1(intermediate_reg_2[77]),.i2(intermediate_reg_2[76]),.o(intermediate_reg_3[38])); 
xor_module xor_module_inst_3_64(.clk(clk),.reset(reset),.i1(intermediate_reg_2[75]),.i2(intermediate_reg_2[74]),.o(intermediate_reg_3[37])); 
mux_module mux_module_inst_3_65(.clk(clk),.reset(reset),.i1(intermediate_reg_2[73]),.i2(intermediate_reg_2[72]),.o(intermediate_reg_3[36]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_66(.clk(clk),.reset(reset),.i1(intermediate_reg_2[71]),.i2(intermediate_reg_2[70]),.o(intermediate_reg_3[35]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_67(.clk(clk),.reset(reset),.i1(intermediate_reg_2[69]),.i2(intermediate_reg_2[68]),.o(intermediate_reg_3[34]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_68(.clk(clk),.reset(reset),.i1(intermediate_reg_2[67]),.i2(intermediate_reg_2[66]),.o(intermediate_reg_3[33])); 
xor_module xor_module_inst_3_69(.clk(clk),.reset(reset),.i1(intermediate_reg_2[65]),.i2(intermediate_reg_2[64]),.o(intermediate_reg_3[32])); 
xor_module xor_module_inst_3_70(.clk(clk),.reset(reset),.i1(intermediate_reg_2[63]),.i2(intermediate_reg_2[62]),.o(intermediate_reg_3[31])); 
xor_module xor_module_inst_3_71(.clk(clk),.reset(reset),.i1(intermediate_reg_2[61]),.i2(intermediate_reg_2[60]),.o(intermediate_reg_3[30])); 
mux_module mux_module_inst_3_72(.clk(clk),.reset(reset),.i1(intermediate_reg_2[59]),.i2(intermediate_reg_2[58]),.o(intermediate_reg_3[29]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_73(.clk(clk),.reset(reset),.i1(intermediate_reg_2[57]),.i2(intermediate_reg_2[56]),.o(intermediate_reg_3[28]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_74(.clk(clk),.reset(reset),.i1(intermediate_reg_2[55]),.i2(intermediate_reg_2[54]),.o(intermediate_reg_3[27]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_75(.clk(clk),.reset(reset),.i1(intermediate_reg_2[53]),.i2(intermediate_reg_2[52]),.o(intermediate_reg_3[26])); 
xor_module xor_module_inst_3_76(.clk(clk),.reset(reset),.i1(intermediate_reg_2[51]),.i2(intermediate_reg_2[50]),.o(intermediate_reg_3[25])); 
mux_module mux_module_inst_3_77(.clk(clk),.reset(reset),.i1(intermediate_reg_2[49]),.i2(intermediate_reg_2[48]),.o(intermediate_reg_3[24]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_78(.clk(clk),.reset(reset),.i1(intermediate_reg_2[47]),.i2(intermediate_reg_2[46]),.o(intermediate_reg_3[23]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_79(.clk(clk),.reset(reset),.i1(intermediate_reg_2[45]),.i2(intermediate_reg_2[44]),.o(intermediate_reg_3[22]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_80(.clk(clk),.reset(reset),.i1(intermediate_reg_2[43]),.i2(intermediate_reg_2[42]),.o(intermediate_reg_3[21])); 
mux_module mux_module_inst_3_81(.clk(clk),.reset(reset),.i1(intermediate_reg_2[41]),.i2(intermediate_reg_2[40]),.o(intermediate_reg_3[20]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_82(.clk(clk),.reset(reset),.i1(intermediate_reg_2[39]),.i2(intermediate_reg_2[38]),.o(intermediate_reg_3[19])); 
xor_module xor_module_inst_3_83(.clk(clk),.reset(reset),.i1(intermediate_reg_2[37]),.i2(intermediate_reg_2[36]),.o(intermediate_reg_3[18])); 
mux_module mux_module_inst_3_84(.clk(clk),.reset(reset),.i1(intermediate_reg_2[35]),.i2(intermediate_reg_2[34]),.o(intermediate_reg_3[17]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_85(.clk(clk),.reset(reset),.i1(intermediate_reg_2[33]),.i2(intermediate_reg_2[32]),.o(intermediate_reg_3[16]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_86(.clk(clk),.reset(reset),.i1(intermediate_reg_2[31]),.i2(intermediate_reg_2[30]),.o(intermediate_reg_3[15])); 
mux_module mux_module_inst_3_87(.clk(clk),.reset(reset),.i1(intermediate_reg_2[29]),.i2(intermediate_reg_2[28]),.o(intermediate_reg_3[14]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_88(.clk(clk),.reset(reset),.i1(intermediate_reg_2[27]),.i2(intermediate_reg_2[26]),.o(intermediate_reg_3[13])); 
xor_module xor_module_inst_3_89(.clk(clk),.reset(reset),.i1(intermediate_reg_2[25]),.i2(intermediate_reg_2[24]),.o(intermediate_reg_3[12])); 
xor_module xor_module_inst_3_90(.clk(clk),.reset(reset),.i1(intermediate_reg_2[23]),.i2(intermediate_reg_2[22]),.o(intermediate_reg_3[11])); 
mux_module mux_module_inst_3_91(.clk(clk),.reset(reset),.i1(intermediate_reg_2[21]),.i2(intermediate_reg_2[20]),.o(intermediate_reg_3[10]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_92(.clk(clk),.reset(reset),.i1(intermediate_reg_2[19]),.i2(intermediate_reg_2[18]),.o(intermediate_reg_3[9]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_93(.clk(clk),.reset(reset),.i1(intermediate_reg_2[17]),.i2(intermediate_reg_2[16]),.o(intermediate_reg_3[8]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_94(.clk(clk),.reset(reset),.i1(intermediate_reg_2[15]),.i2(intermediate_reg_2[14]),.o(intermediate_reg_3[7]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_95(.clk(clk),.reset(reset),.i1(intermediate_reg_2[13]),.i2(intermediate_reg_2[12]),.o(intermediate_reg_3[6]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_96(.clk(clk),.reset(reset),.i1(intermediate_reg_2[11]),.i2(intermediate_reg_2[10]),.o(intermediate_reg_3[5]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_97(.clk(clk),.reset(reset),.i1(intermediate_reg_2[9]),.i2(intermediate_reg_2[8]),.o(intermediate_reg_3[4])); 
mux_module mux_module_inst_3_98(.clk(clk),.reset(reset),.i1(intermediate_reg_2[7]),.i2(intermediate_reg_2[6]),.o(intermediate_reg_3[3]),.sel(intermediate_reg_2[0])); 
xor_module xor_module_inst_3_99(.clk(clk),.reset(reset),.i1(intermediate_reg_2[5]),.i2(intermediate_reg_2[4]),.o(intermediate_reg_3[2])); 
mux_module mux_module_inst_3_100(.clk(clk),.reset(reset),.i1(intermediate_reg_2[3]),.i2(intermediate_reg_2[2]),.o(intermediate_reg_3[1]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_101(.clk(clk),.reset(reset),.i1(intermediate_reg_2[1]),.i2(intermediate_reg_2[0]),.o(intermediate_reg_3[0]),.sel(intermediate_reg_2[0])); 
always@(posedge clk) begin 
outp [101:0] <= intermediate_reg_3; 
outp[103:102] <= intermediate_reg_3[1:0] ; 
end 
endmodule 
 

module spram_2048_40bit_module_4(input clk, input reset, input[207:0] inp, output reg [159:0] outp); 

spram_2048_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[51:0]),.outp(outp[39:0])); 

spram_2048_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[103:52]),.outp(outp[79:40])); 

spram_2048_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[155:104]),.outp(outp[119:80])); 

spram_2048_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[207:156]),.outp(outp[159:120])); 

endmodule 

module tensor_block_bf16_module_3(input clk, input reset, input[794:0] inp, output reg [815:0] outp); 

tensor_block_bf16_module inst_0 (.clk(clk),.reset(reset),.inp(inp[264:0]),.outp(outp[271:0])); 

tensor_block_bf16_module inst_1 (.clk(clk),.reset(reset),.inp(inp[529:265]),.outp(outp[543:272])); 

tensor_block_bf16_module inst_2 (.clk(clk),.reset(reset),.inp(inp[794:530]),.outp(outp[815:544])); 

endmodule 

module systolic_array_4_fp16bit_1(input clk, input reset, input[417:0] inp, output reg [223:0] outp); 

systolic_array_4_fp16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[417:0]),.outp(outp[223:0])); 

endmodule 

module systolic_array_4_fp16bit_2(input clk, input reset, input[835:0] inp, output reg [447:0] outp); 

systolic_array_4_fp16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[417:0]),.outp(outp[223:0])); 

systolic_array_4_fp16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[835:418]),.outp(outp[447:224])); 

endmodule 


module spram_4096_60bit_module_12(input clk, input reset, input[875:0] inp, output reg [719:0] outp); 

spram_4096_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[72:0]),.outp(outp[59:0])); 

spram_4096_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[145:73]),.outp(outp[119:60])); 

spram_4096_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[218:146]),.outp(outp[179:120])); 

spram_4096_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[291:219]),.outp(outp[239:180])); 

spram_4096_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[364:292]),.outp(outp[299:240])); 

spram_4096_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[437:365]),.outp(outp[359:300])); 

spram_4096_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[510:438]),.outp(outp[419:360])); 

spram_4096_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[583:511]),.outp(outp[479:420])); 

spram_4096_60bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[656:584]),.outp(outp[539:480])); 

spram_4096_60bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[729:657]),.outp(outp[599:540])); 

spram_4096_60bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[802:730]),.outp(outp[659:600])); 

spram_4096_60bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[875:803]),.outp(outp[719:660])); 

endmodule 

module adder_tree_4_8bit_12(input clk, input reset, input[1535:0] inp, output reg [191:0] outp); 

adder_tree_4_8bit inst_0 (.clk(clk),.reset(reset),.inp(inp[127:0]),.outp(outp[15:0])); 

adder_tree_4_8bit inst_1 (.clk(clk),.reset(reset),.inp(inp[255:128]),.outp(outp[31:16])); 

adder_tree_4_8bit inst_2 (.clk(clk),.reset(reset),.inp(inp[383:256]),.outp(outp[47:32])); 

adder_tree_4_8bit inst_3 (.clk(clk),.reset(reset),.inp(inp[511:384]),.outp(outp[63:48])); 

adder_tree_4_8bit inst_4 (.clk(clk),.reset(reset),.inp(inp[639:512]),.outp(outp[79:64])); 

adder_tree_4_8bit inst_5 (.clk(clk),.reset(reset),.inp(inp[767:640]),.outp(outp[95:80])); 

adder_tree_4_8bit inst_6 (.clk(clk),.reset(reset),.inp(inp[895:768]),.outp(outp[111:96])); 

adder_tree_4_8bit inst_7 (.clk(clk),.reset(reset),.inp(inp[1023:896]),.outp(outp[127:112])); 

adder_tree_4_8bit inst_8 (.clk(clk),.reset(reset),.inp(inp[1151:1024]),.outp(outp[143:128])); 

adder_tree_4_8bit inst_9 (.clk(clk),.reset(reset),.inp(inp[1279:1152]),.outp(outp[159:144])); 

adder_tree_4_8bit inst_10 (.clk(clk),.reset(reset),.inp(inp[1407:1280]),.outp(outp[175:160])); 

adder_tree_4_8bit inst_11 (.clk(clk),.reset(reset),.inp(inp[1535:1408]),.outp(outp[191:176])); 

endmodule 

module spram_4096_40bit_module_60(input clk, input reset, input[3179:0] inp, output reg [2399:0] outp); 

spram_4096_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[52:0]),.outp(outp[39:0])); 

spram_4096_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[105:53]),.outp(outp[79:40])); 

spram_4096_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[158:106]),.outp(outp[119:80])); 

spram_4096_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[211:159]),.outp(outp[159:120])); 

spram_4096_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[264:212]),.outp(outp[199:160])); 

spram_4096_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[317:265]),.outp(outp[239:200])); 

spram_4096_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[370:318]),.outp(outp[279:240])); 

spram_4096_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[423:371]),.outp(outp[319:280])); 

spram_4096_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[476:424]),.outp(outp[359:320])); 

spram_4096_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[529:477]),.outp(outp[399:360])); 

spram_4096_40bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[582:530]),.outp(outp[439:400])); 

spram_4096_40bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[635:583]),.outp(outp[479:440])); 

spram_4096_40bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[688:636]),.outp(outp[519:480])); 

spram_4096_40bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[741:689]),.outp(outp[559:520])); 

spram_4096_40bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[794:742]),.outp(outp[599:560])); 

spram_4096_40bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[847:795]),.outp(outp[639:600])); 

spram_4096_40bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[900:848]),.outp(outp[679:640])); 

spram_4096_40bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[953:901]),.outp(outp[719:680])); 

spram_4096_40bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[1006:954]),.outp(outp[759:720])); 

spram_4096_40bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[1059:1007]),.outp(outp[799:760])); 

spram_4096_40bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[1112:1060]),.outp(outp[839:800])); 

spram_4096_40bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[1165:1113]),.outp(outp[879:840])); 

spram_4096_40bit_module inst_22 (.clk(clk),.reset(reset),.inp(inp[1218:1166]),.outp(outp[919:880])); 

spram_4096_40bit_module inst_23 (.clk(clk),.reset(reset),.inp(inp[1271:1219]),.outp(outp[959:920])); 

spram_4096_40bit_module inst_24 (.clk(clk),.reset(reset),.inp(inp[1324:1272]),.outp(outp[999:960])); 

spram_4096_40bit_module inst_25 (.clk(clk),.reset(reset),.inp(inp[1377:1325]),.outp(outp[1039:1000])); 

spram_4096_40bit_module inst_26 (.clk(clk),.reset(reset),.inp(inp[1430:1378]),.outp(outp[1079:1040])); 

spram_4096_40bit_module inst_27 (.clk(clk),.reset(reset),.inp(inp[1483:1431]),.outp(outp[1119:1080])); 

spram_4096_40bit_module inst_28 (.clk(clk),.reset(reset),.inp(inp[1536:1484]),.outp(outp[1159:1120])); 

spram_4096_40bit_module inst_29 (.clk(clk),.reset(reset),.inp(inp[1589:1537]),.outp(outp[1199:1160])); 

spram_4096_40bit_module inst_30 (.clk(clk),.reset(reset),.inp(inp[1642:1590]),.outp(outp[1239:1200])); 

spram_4096_40bit_module inst_31 (.clk(clk),.reset(reset),.inp(inp[1695:1643]),.outp(outp[1279:1240])); 

spram_4096_40bit_module inst_32 (.clk(clk),.reset(reset),.inp(inp[1748:1696]),.outp(outp[1319:1280])); 

spram_4096_40bit_module inst_33 (.clk(clk),.reset(reset),.inp(inp[1801:1749]),.outp(outp[1359:1320])); 

spram_4096_40bit_module inst_34 (.clk(clk),.reset(reset),.inp(inp[1854:1802]),.outp(outp[1399:1360])); 

spram_4096_40bit_module inst_35 (.clk(clk),.reset(reset),.inp(inp[1907:1855]),.outp(outp[1439:1400])); 

spram_4096_40bit_module inst_36 (.clk(clk),.reset(reset),.inp(inp[1960:1908]),.outp(outp[1479:1440])); 

spram_4096_40bit_module inst_37 (.clk(clk),.reset(reset),.inp(inp[2013:1961]),.outp(outp[1519:1480])); 

spram_4096_40bit_module inst_38 (.clk(clk),.reset(reset),.inp(inp[2066:2014]),.outp(outp[1559:1520])); 

spram_4096_40bit_module inst_39 (.clk(clk),.reset(reset),.inp(inp[2119:2067]),.outp(outp[1599:1560])); 

spram_4096_40bit_module inst_40 (.clk(clk),.reset(reset),.inp(inp[2172:2120]),.outp(outp[1639:1600])); 

spram_4096_40bit_module inst_41 (.clk(clk),.reset(reset),.inp(inp[2225:2173]),.outp(outp[1679:1640])); 

spram_4096_40bit_module inst_42 (.clk(clk),.reset(reset),.inp(inp[2278:2226]),.outp(outp[1719:1680])); 

spram_4096_40bit_module inst_43 (.clk(clk),.reset(reset),.inp(inp[2331:2279]),.outp(outp[1759:1720])); 

spram_4096_40bit_module inst_44 (.clk(clk),.reset(reset),.inp(inp[2384:2332]),.outp(outp[1799:1760])); 

spram_4096_40bit_module inst_45 (.clk(clk),.reset(reset),.inp(inp[2437:2385]),.outp(outp[1839:1800])); 

spram_4096_40bit_module inst_46 (.clk(clk),.reset(reset),.inp(inp[2490:2438]),.outp(outp[1879:1840])); 

spram_4096_40bit_module inst_47 (.clk(clk),.reset(reset),.inp(inp[2543:2491]),.outp(outp[1919:1880])); 

spram_4096_40bit_module inst_48 (.clk(clk),.reset(reset),.inp(inp[2596:2544]),.outp(outp[1959:1920])); 

spram_4096_40bit_module inst_49 (.clk(clk),.reset(reset),.inp(inp[2649:2597]),.outp(outp[1999:1960])); 

spram_4096_40bit_module inst_50 (.clk(clk),.reset(reset),.inp(inp[2702:2650]),.outp(outp[2039:2000])); 

spram_4096_40bit_module inst_51 (.clk(clk),.reset(reset),.inp(inp[2755:2703]),.outp(outp[2079:2040])); 

spram_4096_40bit_module inst_52 (.clk(clk),.reset(reset),.inp(inp[2808:2756]),.outp(outp[2119:2080])); 

spram_4096_40bit_module inst_53 (.clk(clk),.reset(reset),.inp(inp[2861:2809]),.outp(outp[2159:2120])); 

spram_4096_40bit_module inst_54 (.clk(clk),.reset(reset),.inp(inp[2914:2862]),.outp(outp[2199:2160])); 

spram_4096_40bit_module inst_55 (.clk(clk),.reset(reset),.inp(inp[2967:2915]),.outp(outp[2239:2200])); 

spram_4096_40bit_module inst_56 (.clk(clk),.reset(reset),.inp(inp[3020:2968]),.outp(outp[2279:2240])); 

spram_4096_40bit_module inst_57 (.clk(clk),.reset(reset),.inp(inp[3073:3021]),.outp(outp[2319:2280])); 

spram_4096_40bit_module inst_58 (.clk(clk),.reset(reset),.inp(inp[3126:3074]),.outp(outp[2359:2320])); 

spram_4096_40bit_module inst_59 (.clk(clk),.reset(reset),.inp(inp[3179:3127]),.outp(outp[2399:2360])); 

endmodule 

module tensor_block_bf16_module_2(input clk, input reset, input[529:0] inp, output reg [543:0] outp); 

tensor_block_bf16_module inst_0 (.clk(clk),.reset(reset),.inp(inp[264:0]),.outp(outp[271:0])); 

tensor_block_bf16_module inst_1 (.clk(clk),.reset(reset),.inp(inp[529:265]),.outp(outp[543:272])); 

endmodule 


module adder_tree_3_fp16bit_8(input clk, input reset, input[1055:0] inp, output reg [127:0] outp); 

adder_tree_3_fp16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[131:0]),.outp(outp[15:0])); 

adder_tree_3_fp16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[263:132]),.outp(outp[31:16])); 

adder_tree_3_fp16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[395:264]),.outp(outp[47:32])); 

adder_tree_3_fp16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[527:396]),.outp(outp[63:48])); 

adder_tree_3_fp16bit inst_4 (.clk(clk),.reset(reset),.inp(inp[659:528]),.outp(outp[79:64])); 

adder_tree_3_fp16bit inst_5 (.clk(clk),.reset(reset),.inp(inp[791:660]),.outp(outp[95:80])); 

adder_tree_3_fp16bit inst_6 (.clk(clk),.reset(reset),.inp(inp[923:792]),.outp(outp[111:96])); 

adder_tree_3_fp16bit inst_7 (.clk(clk),.reset(reset),.inp(inp[1055:924]),.outp(outp[127:112])); 

endmodule 

module spram_2048_40bit_module_2(input clk, input reset, input[103:0] inp, output reg [79:0] outp); 

spram_2048_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[51:0]),.outp(outp[39:0])); 

spram_2048_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[103:52]),.outp(outp[79:40])); 

endmodule 

module adder_tree_3_16bit_4(input clk, input reset, input[511:0] inp, output reg [127:0] outp); 

adder_tree_3_16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[127:0]),.outp(outp[31:0])); 

adder_tree_3_16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[255:128]),.outp(outp[63:32])); 

adder_tree_3_16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[383:256]),.outp(outp[95:64])); 

adder_tree_3_16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[511:384]),.outp(outp[127:96])); 

endmodule 

module adder_tree_3_fp16bit_10(input clk, input reset, input[1319:0] inp, output reg [159:0] outp); 

adder_tree_3_fp16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[131:0]),.outp(outp[15:0])); 

adder_tree_3_fp16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[263:132]),.outp(outp[31:16])); 

adder_tree_3_fp16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[395:264]),.outp(outp[47:32])); 

adder_tree_3_fp16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[527:396]),.outp(outp[63:48])); 

adder_tree_3_fp16bit inst_4 (.clk(clk),.reset(reset),.inp(inp[659:528]),.outp(outp[79:64])); 

adder_tree_3_fp16bit inst_5 (.clk(clk),.reset(reset),.inp(inp[791:660]),.outp(outp[95:80])); 

adder_tree_3_fp16bit inst_6 (.clk(clk),.reset(reset),.inp(inp[923:792]),.outp(outp[111:96])); 

adder_tree_3_fp16bit inst_7 (.clk(clk),.reset(reset),.inp(inp[1055:924]),.outp(outp[127:112])); 

adder_tree_3_fp16bit inst_8 (.clk(clk),.reset(reset),.inp(inp[1187:1056]),.outp(outp[143:128])); 

adder_tree_3_fp16bit inst_9 (.clk(clk),.reset(reset),.inp(inp[1319:1188]),.outp(outp[159:144])); 

endmodule 


module systolic_array_4_fp16bit_3(input clk, input reset, input[1253:0] inp, output reg [671:0] outp); 

systolic_array_4_fp16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[417:0]),.outp(outp[223:0])); 

systolic_array_4_fp16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[835:418]),.outp(outp[447:224])); 

systolic_array_4_fp16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[1253:836]),.outp(outp[671:448])); 

endmodule 


module spram_4096_40bit_module_24(input clk, input reset, input[1271:0] inp, output reg [959:0] outp); 

spram_4096_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[52:0]),.outp(outp[39:0])); 

spram_4096_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[105:53]),.outp(outp[79:40])); 

spram_4096_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[158:106]),.outp(outp[119:80])); 

spram_4096_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[211:159]),.outp(outp[159:120])); 

spram_4096_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[264:212]),.outp(outp[199:160])); 

spram_4096_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[317:265]),.outp(outp[239:200])); 

spram_4096_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[370:318]),.outp(outp[279:240])); 

spram_4096_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[423:371]),.outp(outp[319:280])); 

spram_4096_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[476:424]),.outp(outp[359:320])); 

spram_4096_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[529:477]),.outp(outp[399:360])); 

spram_4096_40bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[582:530]),.outp(outp[439:400])); 

spram_4096_40bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[635:583]),.outp(outp[479:440])); 

spram_4096_40bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[688:636]),.outp(outp[519:480])); 

spram_4096_40bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[741:689]),.outp(outp[559:520])); 

spram_4096_40bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[794:742]),.outp(outp[599:560])); 

spram_4096_40bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[847:795]),.outp(outp[639:600])); 

spram_4096_40bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[900:848]),.outp(outp[679:640])); 

spram_4096_40bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[953:901]),.outp(outp[719:680])); 

spram_4096_40bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[1006:954]),.outp(outp[759:720])); 

spram_4096_40bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[1059:1007]),.outp(outp[799:760])); 

spram_4096_40bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[1112:1060]),.outp(outp[839:800])); 

spram_4096_40bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[1165:1113]),.outp(outp[879:840])); 

spram_4096_40bit_module inst_22 (.clk(clk),.reset(reset),.inp(inp[1218:1166]),.outp(outp[919:880])); 

spram_4096_40bit_module inst_23 (.clk(clk),.reset(reset),.inp(inp[1271:1219]),.outp(outp[959:920])); 

endmodule 


module adder_tree_1_16bit (input clk,input reset,input [31:0] inp, output reg [31:0] outp);

adder_tree_1stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.sum_out(outp));

endmodule

module adder_tree_2_16bit (input clk, input reset, input [63:0] inp, output reg [31:0] outp);

adder_tree_2stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.sum_out(outp));

endmodule

module adder_tree_3_16bit (input clk, input reset, input [127:0] inp, output reg [31:0] outp);

adder_tree_3stage_16bit inst (.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.inp20(inp[79:64]),.inp21(inp[95:80]),.inp30(inp[111:96]),.inp31(inp[127:112]),.sum_out(outp));

endmodule

module adder_tree_4_16bit (input clk, input reset, input [255:0] inp, output reg [31:0] outp);

adder_tree_4stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.inp20(inp[79:64]),.inp21(inp[95:80]),.inp30(inp[111:96]),.inp31(inp[127:112]),.inp40(inp[143:128]),.inp41(inp[159:144]),.inp50(inp[175:160]),.inp51(inp[191:176]),.inp60(inp[207:192]),.inp61(inp[223:208]),.inp70(inp[239:224]),.inp71(inp[255:240]),.sum_out(outp));

endmodule

module adder_tree_1_8bit (input clk, input reset, input [15:0] inp, output reg [15:0] outp);

adder_tree_1stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.sum_out(outp));

endmodule

module adder_tree_2_8bit (input clk, input reset, input [31:0] inp, output reg [15:0] outp);

adder_tree_2stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.sum_out(outp));

endmodule

module adder_tree_3_8bit (input clk, input reset, input [63:0] inp, output reg [15:0] outp);

adder_tree_3stage_8bit inst (.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.inp20(inp[39:32]),.inp21(inp[47:40]),.inp30(inp[55:48]),.inp31(inp[63:56]),.sum_out(outp));

endmodule

module adder_tree_4_8bit (input clk, input reset, input [127:0] inp, output reg [15:0] outp);

adder_tree_4stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.inp20(inp[39:32]),.inp21(inp[47:40]),.inp30(inp[55:48]),.inp31(inp[63:56]),.inp40(inp[71:64]),.inp41(inp[79:72]),.inp50(inp[87:80]),.inp51(inp[95:88]),.inp60(inp[103:96]),.inp61(inp[111:104]),.inp70(inp[119:112]),.inp71(inp[127:120]),.sum_out(outp));

endmodule

module adder_tree_1_4bit (input clk, input reset, input [7:0] inp, output reg [7:0] outp);

adder_tree_1stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.sum_out(outp));

endmodule

module adder_tree_2_4bit (input clk, input reset, input [15:0] inp, output reg [7:0] outp);

adder_tree_2stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.sum_out(outp));

endmodule

module adder_tree_3_4bit (input clk, input reset, input [31:0] inp, output reg [7:0] outp);

adder_tree_3stage_4bit inst (.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.inp20(inp[19:16]),.inp21(inp[23:20]),.inp30(inp[27:24]),.inp31(inp[31:28]),.sum_out(outp));

endmodule

module adder_tree_4_4bit (input clk, input reset, input [63:0] inp, output reg [7:0] outp);

adder_tree_4stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.inp20(inp[19:16]),.inp21(inp[23:20]),.inp30(inp[27:24]),.inp31(inp[31:28]),.inp40(inp[35:32]),.inp41(inp[39:36]),.inp50(inp[43:40]),.inp51(inp[47:44]),.inp60(inp[51:48]),.inp61(inp[55:52]),.inp70(inp[59:56]),.inp71(inp[63:60]),.sum_out(outp));

endmodule

module adder_tree_3_fp16bit (input clk, input reset, input [131:0] inp, output reg [15:0] outp);

mode4_adder_tree inst(
  .inp0(inp[15:0]),
  .inp1(inp[31:16]),
  .inp2(inp[47:32]),
  .inp3(inp[63:48]),
  .inp4(inp[79:64]),
  .inp5(inp[95:80]),
  .inp6(inp[111:96]),
  .inp7(inp[127:112]),
  .mode4_stage0_run(inp[128]),
  .mode4_stage1_run(inp[129]),
  .mode4_stage2_run(inp[130]),
  .mode4_stage3_run(inp[131]),

  .clk(clk),
  .reset(reset),
  .outp(outp[15:0])
);

endmodule

module dpram_1024_32bit_module (input clk, input reset, input [85:0] inp, output reg [63:0] outp);

dpram inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[53:22]),.data_b(inp[85:54]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_1024_64bit_module (input clk, input reset, input [149:0] inp, output reg [63:0] outp );

dpram_1024_64bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[85:22]),.data_b(inp[149:86]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_2048_64bit_module (input clk, input reset, input [151:0] inp, output reg [127:0] outp);

dpram_2048_64bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[87:24]),.data_b(inp[151:88]),.out_a(outp[63:0]),.out_b(outp[127:64]));

endmodule

module dpram_2048_32bit_module (input clk, input reset, input [87:0] inp, output reg [63:0] outp);

dpram_2048_32bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[55:24]),.data_b(inp[87:56]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_1024_40bit_module (input clk, input reset, input [101:0] inp, output reg [79:0] outp);

dpram_1024_40bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[61:22]),.data_b(inp[101:62]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_1024_60bit_module (input clk, input reset, input [141:0] inp, output reg [119:0] outp);

dpram_1024_60bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[81:22]),.data_b(inp[141:82]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dpram_2048_40bit_module (input clk, input reset, input [103:0] inp, output reg [79:0] outp);

dpram_2048_40bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[63:24]),.data_b(inp[103:64]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_2048_60bit_module (input clk, input reset, input [143:0] inp, output reg [119:0] outp);

dpram_2048_60bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[83:24]),.data_b(inp[143:84]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dpram_4096_40bit_module (input clk, input reset, input [105:0] inp, output reg [79:0] outp);

dpram_4096_40bit inst (.clk(clk),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[65:26]),.data_b(inp[105:66]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_4096_60bit_module (input clk, input reset, input [145:0] inp, output reg [119:0] outp);

dpram_4096_60bit inst (.clk(clk),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[85:26]),.data_b(inp[145:86]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module spram_1024_32bit_module (input clk,input reset,input [42:0] inp, output reg [31:0] outp);

spram inst (.clk(clk),.address(inp[9:0]),.wren(inp[10]),.data(inp[42:11]),.out(outp));

endmodule

module spram_2048_40bit_module (input clk,input reset,input [51:0] inp, output reg [39:0] outp);

spram_2048_40bit inst (.clk(clk),.address(inp[10:0]),.wren(inp[11]),.data(inp[51:12]),.out(outp));

endmodule

module spram_2048_60bit_module (input clk,input reset,input [71:0] inp, output reg [59:0] outp);

spram_2048_60bit inst (.clk(clk),.address(inp[10:0]),.wren(inp[11]),.data(inp[71:12]),.out(outp));

endmodule

module spram_4096_40bit_module (input clk,input reset,input [52:0] inp, output reg [39:0] outp);

spram_4096_40bit inst (.clk(clk),.address(inp[11:0]),.wren(inp[12]),.data(inp[52:13]),.out(outp));

endmodule

module spram_4096_60bit_module (input clk,input reset,input [72:0] inp, output reg [59:0] outp);

spram_4096_60bit inst (.clk(clk),.address(inp[11:0]),.wren(inp[12]),.data(inp[72:13]),.out(outp));

endmodule

module dbram_2048_40bit_module (input clk,input reset,input [103:0] inp, output reg [79:0] outp);

dbram_2048_40bit inst (.clk(clk),.reset(reset),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[63:24]),.data_b(inp[103:64]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dbram_2048_60bit_module (input clk,input reset,input [143:0] inp, output reg [119:0] outp);

dbram_2048_60bit inst (.clk(clk),.reset(reset),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[83:24]),.data_b(inp[143:84]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dbram_4096_40bit_module (input clk,input reset,input [105:0] inp, output reg [79:0] outp);

dbram_4096_40bit inst (.clk(clk),.reset(reset),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[65:26]),.data_b(inp[105:66]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dbram_4096_60bit_module (input clk,input reset,input [145:0] inp, output reg [119:0] outp);

dbram_4096_60bit inst (.clk(clk),.reset(reset),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[85:26]),.data_b(inp[145:86]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule


module fifo_256_40bit_module (input clk,input reset,input [42:0] inp, output reg [41:0] outp);

fifo_256_40bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[40:1]),.we(inp[41]),.dout(outp[39:0]),.re(inp[42]),.full(outp[40]),.empty(outp[41]));

endmodule

module fifo_256_60bit_module (input clk,input reset,input [62:0] inp, output reg [61:0] outp);

fifo_256_60bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[60:1]),.we(inp[61]),.dout(outp[59:0]),.re(inp[62]),.full(outp[60]),.empty(outp[61]));

endmodule

module fifo_512_60bit_module (input clk,input reset,input [62:0] inp, output reg [61:0] outp);

fifo_512_60bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[60:1]),.we(inp[61]),.dout(outp[59:0]),.re(inp[62]),.full(outp[60]),.empty(outp[61]));

endmodule

module fifo_512_40bit_module (input clk,input reset,input [42:0] inp, output reg [41:0] outp);

fifo_512_40bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[40:1]),.we(inp[41]),.dout(outp[39:0]),.re(inp[42]),.full(outp[40]),.empty(outp[41]));

endmodule

module tanh_16bit (input clk,input reset, input [15:0] inp, output reg [15:0] outp);

tanh inst (.x(inp),.tanh_out(outp));

endmodule

module sigmoid_16bit (input clk,input reset, input [15:0] inp, output reg [15:0] outp);

sigmoid inst (.x(inp),.sig_out(outp));

endmodule

module systolic_array_4_16bit (input clk, input reset, input [254:0] inp, output reg [130:0] outp);

matmul_4x4_systolic inst(
 .clk(clk),
 .reset(inp[254]),
 .pe_reset(reset),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[11:1]),
 .address_mat_b(inp[22:12]),
 .address_mat_c(inp[33:23]),
 .address_stride_a(inp[41:34]),
 .address_stride_b(inp[49:42]),
 .address_stride_c(inp[57:50]),
 .a_data(inp[89:58]),
 .b_data(inp[121:90]),
 .a_data_in(inp[153:122]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[185:154]),
 .c_data_in(inp[217:186]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[32:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[64:33]),
 .b_data_out(outp[96:65]),
 .a_addr(outp[107:97]),
 .b_addr(outp[118:108]),
 .c_addr(outp[129:119]),
 .c_data_available(outp[130]),
 .validity_mask_a_rows(inp[221:218]),
 .validity_mask_a_cols_b_rows(inp[225:222]),
 .validity_mask_b_cols(inp[229:226]),
 .final_mat_mul_size(inp[237:230]),
 .a_loc(inp[245:238]),
 .b_loc(inp[253:246])
);

endmodule

module systolic_array_8_16bit (input clk, input reset, input [785:0] inp, output reg [433:0] outp);

matmul_8x8_systolic inst(
 .clk(clk),
 .reset(reset),
 .pe_reset(inp[785]),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[16:1]),
 .address_mat_b(inp[32:17]),
 .address_mat_c(inp[48:33]),
 .address_stride_a(inp[64:49]),
 .address_stride_b(inp[80:65]),
 .address_stride_c(inp[96:81]),
 .a_data(inp[224:97]),
 .b_data(inp[352:225]),
 .a_data_in(inp[480:353]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[608:481]),
 .c_data_in(inp[736:609]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[128:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[256:129]),
 .b_data_out(outp[384:257]),
 .a_addr(outp[400:385]),
 .b_addr(outp[416:401]),
 .c_addr(outp[432:417]),
 .c_data_available(outp[433]),
 .validity_mask_a_rows(inp[744:737]),
 .validity_mask_a_cols_b_rows(inp[752:745]),
 .validity_mask_b_cols(inp[760:753]),
 .final_mat_mul_size(inp[768:761]),
 .a_loc(inp[776:769]),
 .b_loc(inp[784:777])
);

endmodule

module systolic_array_4_fp16bit (input clk, input reset, input [417:0] inp, output reg [223:0] outp);

matmul_4x4_fp_systolic inst(
 .clk(clk),
 .reset(reset),
 .pe_reset(inp[417]),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[10:1]),
 .address_mat_b(inp[20:11]),
 .address_mat_c(inp[30:21]),
 .address_stride_a(inp[40:31]),
 .address_stride_b(inp[50:41]),
 .address_stride_c(inp[60:51]),
 .a_data(inp[124:61]),
 .b_data(inp[188:125]),
 .a_data_in(inp[252:189]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[316:253]),
 .c_data_in(inp[380:317]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[64:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[128:65]),
 .b_data_out(outp[192:129]),
 .a_addr(outp[202:193]),
 .b_addr(outp[212:203]),
 .c_addr(outp[222:213]),
 .c_data_available(outp[223]),
 .validity_mask_a_rows(inp[384:381]),
 .validity_mask_a_cols_b_rows(inp[388:385]),
 .validity_mask_b_cols(inp[392:389]),
 .final_mat_mul_size(inp[400:393]),
 .a_loc(inp[408:401]),
 .b_loc(inp[416:409])
);

endmodule

module dsp_chain_2_int_sop_2_module (input clk, input reset, input [147:0] inp, output reg [36:0] outp);

dsp_chain_2_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.result(outp[36:0]));

endmodule

module dsp_chain_3_int_sop_2_module (input clk, input reset, input [221:0] inp, output reg [36:0] outp);

dsp_chain_3_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.ax3(inp[165:148]),.ay3(inp[184:166]),.bx3(inp[202:185]),.by3(inp[221:203]),.result(outp[36:0]));

endmodule

module dsp_chain_4_int_sop_2_module (input clk, input reset, input [295:0] inp, output reg [36:0] outp);

dsp_chain_4_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.ax3(inp[165:148]),.ay3(inp[184:166]),.bx3(inp[202:185]),.by3(inp[221:203]),.ax4(inp[239:222]),.ay4(inp[258:240]),.bx4(inp[276:259]),.by4(inp[295:277]),.result(outp[36:0]));

endmodule

module dsp_chain_2_fp16_sop2_mult_module (input clk, input reset, input [127:0] inp, output reg [31:0] outp);

dsp_chain_2_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.result(outp));

endmodule

module dsp_chain_3_fp16_sop2_mult_module (input clk, input reset, input [191:0] inp, output reg [31:0] outp);

dsp_chain_3_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.top_a3(inp[143:128]),.top_b3(inp[159:144]),.bot_a3(inp[175:160]),.bot_b3(inp[191:176]),.result(outp));

endmodule

module dsp_chain_4_fp16_sop2_mult_module (input clk, input reset, input [255:0] inp, output reg [31:0] outp);

dsp_chain_4_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.top_a3(inp[143:128]),.top_b3(inp[159:144]),.bot_a3(inp[175:160]),.bot_b3(inp[191:176]),.top_a4(inp[207:192]),.top_b4(inp[223:208]),.bot_a4(inp[239:224]),.bot_b4(inp[255:240]),.result(outp));

endmodule

module tensor_block_bf16_module (input clk, input reset, input [264:0] inp, output reg [271:0] outp);

tensor_block_bf16 inst(
	.clk(clk),
	.reset(reset),

	.data_in(inp[79:0]),
	.cascade_in(inp[159:80]),
	.acc0_in(inp[191:160]),
	.acc1_in(inp[223:192]),
	.acc2_in(inp[255:224]),
	.accumulator_input1_select(inp[258:256]),

	.out0(outp[31:0]),
	.out1(outp[63:32]),
	.out2(outp[95:64]),
	.cascade_out(outp[175:96]),
	.acc0_out(outp[207:176]),
	.acc1_out(outp[239:208]),
	.acc2_out(outp[271:240]),

	.mux1_select(inp[259]),
	.dot_unit_input_1_enable(inp[260]),
	.bank0_data_in_enable(inp[261]),
	.bank1_data_in_enable(inp[262]),
	.cascade_out_select(inp[263]),
	.dot_unit_input_2_select(inp[264])

	);

endmodule

module tensor_block_int8_module (input clk, input reset, input [264:0] inp, output reg [250:0] outp);

tensor_block inst(
	.clk(clk),
	.reset(reset),

	.data_in(inp[79:0]),
	.cascade_in(inp[159:80]),
	.acc0_in(inp[191:160]),
	.acc1_in(inp[223:192]),
	.acc2_in(inp[255:224]),
	.accumulator_input1_select(inp[258:256]),

	.out0(outp[24:0]),
	.out1(outp[49:25]),
	.out2(outp[74:50]),
	.cascade_out(outp[154:75]),
	.acc0_out(outp[186:155]),
	.acc1_out(outp[218:187]),
	.acc2_out(outp[250:219]),

	.mux1_select(inp[259]),
	.dot_unit_input_1_enable(inp[260]),
	.bank0_data_in_enable(inp[261]),
	.bank1_data_in_enable(inp[262]),
	.cascade_out_select(inp[263]),
	.dot_unit_input_2_select(inp[264])

	);

endmodule


module activation_32_8bit_module (input clk, input reset, input [260:0] inp, output reg [257:0] outp);

activation_32_8bit inst (
    .activation_type(inp[0]),
    .enable_activation(inp[1]),
    .in_data_available(inp[2]),
    .inp_data(inp[258:3]),
    .out_data(outp[255:0]),
    .out_data_available(outp[256]),
    .validity_mask(inp[260:259]),
    .done_activation(outp[257]),
    .clk(clk),
    .reset(reset)
);

endmodule

module activation_32_16bit_module (input clk, input reset, input [515:0] inp, output reg [513:0] outp);

activation_32_16bit inst (
    .activation_type(inp[0]),
    .enable_activation(inp[1]),
    .in_data_available(inp[2]),
    .inp_data(inp[514:3]),
    .out_data(outp[511:0]),
    .out_data_available(outp[512]),
    .validity_mask(inp[515:514]),
    .done_activation(outp[513]),
    .clk(clk),
    .reset(reset)
);

endmodule

module fsm(input clk, input reset, input i1, input i2, output reg o);
// mealy machine

reg [1:0] current_state; 
reg [1:0] next_state;

wire [1:0] inp; 
assign inp = {i2,i1}; 

always@(posedge clk) begin 
	if (reset == 1'b1) begin 
		current_state <= 1'b0; 
	end
	else begin 
		current_state <= next_state; 
	end
end

always@(posedge clk) begin 

	next_state = current_state; 

	case(current_state)
		2'b00:	begin 
							if(inp == 2'b00) begin 
								next_state <= 2'b00; 
								o <= 1'b0; 
							end
							if (inp == 2'b01) begin 
								next_state <= 2'b11;
								o <= 1'b1;
							end
							if(inp == 2'b10) begin
  							next_state <= 2'b01;
  							o <= 1'b0;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b10;
							  o <= 1'b0;
							end
					 	end 
		2'b01:	begin 
							if(inp == 2'b00) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b01;
							  o <= 1'b0;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b00;
							  o <= 1'b1;
							end
						end
		2'b10:	begin 
							if(inp == 2'b00) begin
							  next_state <= 2'b11;
							  o <= 1'b0;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b11;
							  o <= 1'b0;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
						end
		2'b11:	begin 
							if(inp == 2'b00) begin
  							next_state <= 2'b00;
							  o <= 1'b1;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b11;
							  o <= 1'b1;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
						end
//		defualt:	begin  
//								next_state <= 2'b00;
//								o <= 1'b0; 
//							end
	endcase
end 

endmodule 
module xor_module (input clk, input reset, input i1, input i2, output reg o);

always@(posedge clk) begin 
if (reset ==1'b1) begin 
o<= 1'b0; 
end
else begin
o <= i1^i2; 
end 
end
endmodule
module mux_module (input clk, input reset, input i1, input i2, output reg o, input sel);

always@(posedge clk) begin 
if (reset ==1'b1) begin 
	o<= 1'b0; 
end

else begin
	if (sel == 1'b0) begin 
		o <= i1;
	end
	else begin
		o <= i2; 
	end 
end 

end

endmodule

`ifdef complex_dsp
module int_sop_2_dspchain (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
	chainin,
	resulta,
	chainout);
input [10:0] mode_sigs;
input clk;
input reset; 
input [17:0] ax, bx;
input [18:0] ay, by;
input [36:0] chainin;

output reg [36:0] resulta;
output reg [36:0] chainout;

wire [11:0] mode_sigs_int;
assign mode_sigs_int = {1'b0, mode_sigs};

int_sop_2 inst1(.clk(clk),.reset(reset),.ax(ax),.bx(bx),.ay(ay),.by(by),.mode_sigs(mode_sigs_int),.chainin(chainin),.result(resulta),.chainout(chainout)); 

endmodule
`else
module int_sop_2_dspchain (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
	chainin,
	resulta,
	chainout);
input [10:0] mode_sigs;
input clk;
input reset; 
input [17:0] ax, bx;
input [18:0] ay, by;
input [36:0] chainin;

output reg [36:0] resulta;
output reg [36:0] chainout;
reg [17:0] ax_reg;
reg [18:0] ay_reg;
reg [17:0] bx_reg;
reg [18:0] by_reg;
reg [36:0] resulta;
always @(posedge clk) begin
  if(reset) begin
    resulta <= 0;
    ax_reg <= 0;
    ay_reg <= 0;
    bx_reg <= 0;
    by_reg <= 0;
  end
  else begin
    ax_reg <= ax;
    ay_reg <= ay;
    bx_reg <= bx;
    by_reg <= by;
    resulta <= ax_reg * ay_reg + bx_reg * by_reg + chainin;
  end
end
assign chainout = resulta;
endmodule
`endif

`ifdef complex_dsp
module fp16_sop2_mult_dspchain (clk,reset,top_a,top_b,bot_a,bot_b,fp32_in,mode_sigs,chainin,chainout,result);
input clk; 
input reset;
input [10:0] mode_sigs; 
input [15:0] top_a,top_b,bot_a,bot_b;
input [31:0] chainin,fp32_in; 
output reg [31:0] chainout, result;

fp16_sop2_mult inst1(.clk(clk),.reset(reset),.top_a(top_a),.top_b(top_b),.bot_a(bot_a),.bot_b(bot_b),.fp32_in(fp32_in),.mode_sigs(mode_sigs),.chainin(chainin),.chainout(chainout),.result(result)); 

endmodule

`else
module fp16_sop2_mult_dspchain (clk,reset,top_a,top_b,bot_a,bot_b,fp32_in,mode_sigs,chainin,chainout,result);
input clk; 
input reset;
input [10:0] mode_sigs; 
input [15:0] top_a,top_b,bot_a,bot_b;
input [31:0] chainin,fp32_in; 
output reg [31:0] chainout, result; 

reg [15:0] top_a_reg,top_b_reg,bot_a_reg,bot_b_reg; 
reg [31:0] chainin_reg; 
reg [31:0] r1,r2,r3; 
always@(posedge clk) begin 
if(reset) begin 
top_a_reg<= 16'b0; 
top_b_reg<= 16'b0; 
bot_a_reg<= 16'b0; 
bot_b_reg<= 16'b0;
//result<=32'b0;
//chainout<=32'b0;
chainin_reg<=32'b0;   
end
else begin 
top_a_reg<=top_a; 
top_b_reg<=top_b; 
bot_a_reg<=bot_a;
bot_b_reg<=bot_b;
//chainout<=result;
chainin_reg<=chainin; 
end
end

wire [4:0] flags1,flags2,flags3,flags4; 

FPMult_16_dspchain inst1(.clk(clk),.rst(reset),.a(top_a_reg),.b(top_b_reg),.flags(flags1),.result(r1)); 
FPMult_16_dspchain inst2(.clk(clk),.rst(reset),.a(bot_a_reg),.b(bot_b_reg),.flags(flags2),.result(r2));
FPAddSub_single_dspchain inst3(.clk(clk),.rst(reset),.a(r1),.b(r2),.flags(flags3),.operation(1'b1),.result(r3));
FPAddSub_single_dspchain inst4(.clk(clk),.rst(reset),.a(r3),.b(chainin),.flags(flags4),.operation(1'b1),.result(result));
assign chainout = result; 
endmodule
//`endif

//`timescale 1ns / 1ps


// IEEE Half Precision => 5 = 5, 10 = 10



//`define IEEE_COMPLIANCE 1


//////////////////////////////////////////////////////////////////////////////////
//
// Module Name:    FPMult
//
//////////////////////////////////////////////////////////////////////////////////

module FPMult_16_dspchain(
		clk,
		rst,
		a,
		b,
		result,
		flags
    );
	
	// Input Ports
	input clk ;							// Clock
	input rst ;							// Reset signal
	input [16-1:0] a;						// Input A, a 32-bit floating point number
	input [16-1:0] b;						// Input B, a 32-bit floating point number
	
	// Output ports
	output [32-1:0] result ;					// Product, result of the operation, 32-bit FP number
	output [4:0] flags ;						// Flags indicating exceptions according to IEEE754
	
	// Internal signals
	wire [32-1:0] Z_int ;					// Product, result of the operation, 32-bit FP number
	wire [4:0] Flags_int ;						// Flags indicating exceptions according to IEEE754
	
	wire Sa ;							// A's sign
	wire Sb ;							// B's sign
	wire Sp ;							// Product sign
	wire [5-1:0] Ea ;					// A's 5
	wire [5-1:0] Eb ;					// B's 5
	wire [2*10+1:0] Mp ;					// Product 10
	wire [4:0] InputExc ;						// Exceptions in inputs
	wire [23-1:0] NormM ;					// Normalized 10
	wire [8:0] NormE ;					// Normalized 5
	wire [23:0] RoundM ;					// Normalized 10
	wire [8:0] RoundE ;					// Normalized 5
	wire [23:0] RoundMP ;					// Normalized 10
	wire [8:0] RoundEP ;					// Normalized 5
	wire GRS ;

	//reg [63:0] pipe_0;						// Pipeline register Input->Prep
	reg [2*16-1:0] pipe_0;					// Pipeline register Input->Prep

	//reg [92:0] pipe_1;						// Pipeline register Prep->Execute
	//reg [3*10+2*5+7:0] pipe_1;			// Pipeline register Prep->Execute
	reg [3*10+2*5+18:0] pipe_1;

	//reg [38:0] pipe_2;						// Pipeline register Execute->Normalize
	reg [23+8+7:0] pipe_2;				// Pipeline register Execute->Normalize

	//reg [72:0] pipe_3;						// Pipeline register Normalize->Round
	reg [2*23+2*8+10:0] pipe_3;			// Pipeline register Normalize->Round

	//reg [36:0] pipe_4;						// Pipeline register Round->Output
	reg [32+4:0] pipe_4;					// Pipeline register Round->Output
	
	assign result = pipe_4[32+4:5] ;
	assign flags = pipe_4[4:0] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPMult_PrepModule_dspchain PrepModule(clk, rst, pipe_0[2*16-1:16], pipe_0[16-1:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10+1:0], InputExc[4:0]) ;

	// Perform (unsigned) 10 multiplication
	FPMult_ExecuteModule_dspchain ExecuteModule(pipe_1[3*10+5*2+7:2*10+2*5+8], pipe_1[2*10+2*5+7:2*10+7], pipe_1[2*10+6:5], pipe_1[2*10+2*5+6:2*10+5+7], pipe_1[2*10+5+6:2*10+7], pipe_1[2*10+2*5+8], pipe_1[2*10+2*5+7], Sp, NormE[8:0], NormM[23-1:0], GRS) ;

	// Round result and if necessary, perform a second (post-rounding) normalization step
	FPMult_NormalizeModule_dspchain NormalizeModule(pipe_2[23-1:0], pipe_2[23+8:23], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]) ;		

	// Round result and if necessary, perform a second (post-rounding) normalization step
	//FPMult_RoundModule RoundModule(pipe_3[47:24], pipe_3[23:0], pipe_3[65:57], pipe_3[56:48], pipe_3[66], pipe_3[67], pipe_3[72:68], Z_int[31:0], Flags_int[4:0]) ;		
	FPMult_RoundModule_dspchain RoundModule(pipe_3[2*23+1:23+1], pipe_3[23:0], pipe_3[2*8+2*23+3:2*23+8+3], pipe_3[2*23+8+2:2*23+2], pipe_3[2*23+2*8+4], pipe_3[2*23+2*8+5], pipe_3[2*23+2*8+10:2*23+2*8+6], Z_int[32-1:0], Flags_int[4:0]) ;		


//adding always@ (*) instead of posedge clock to make design combinational
	always @ (*) begin	
		if(rst) begin
			pipe_0 = 0;
			pipe_1 = 0;
			pipe_2 = 0; 
			pipe_3 = 0;
			pipe_4 = 0;
		end 
		else begin		
			/* PIPE 0
				[2*16-1:16] A
				[16-1:0] B
			*/
                       pipe_0 = {a, b} ;


			/* PIPE 1
				[2*5+3*10 + 18: 2*5+2*10 + 18] //pipe_0[16+10-1:16] , 10 of A
				[2*5+2*10 + 17 :2*5+2*10 + 9] // pipe_0[8:0]
				[2*5+2*10 + 8] Sa
				[2*5+2*10 + 7] Sb
				[2*5+2*10 + 6:5+2*10+7] Ea
				[5 +2*10+6:2*10+7] Eb
				[2*10+1+5:5] Mp
				[4:0] InputExc
			*/
			//pipe_1 <= {pipe_0[16+10-1:16], pipe_0[10_MUL_SPLIT_LSB-1:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10-1:0], InputExc[4:0]} ;
			pipe_1 = {pipe_0[16+10-1:16], pipe_0[8:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10+1:0], InputExc[4:0]} ;
			
			/* PIPE 2
				[8 + 23 + 7:8 + 23 + 3] InputExc
				[8 + 23 + 2] GRS
				[8 + 23 + 1] Sp
				[8 + 23:23] NormE
				[23-1:0] NormM
			*/
			pipe_2 = {pipe_1[4:0], GRS, Sp, NormE[8:0], NormM[23-1:0]} ;
			/* PIPE 3
				[2*8+2*23+10:2*8+2*23+6] InputExc
				[2*8+2*23+5] GRS
				[2*8+2*23+4] Sp	
				[2*8+2*23+3:8+2*23+3] RoundE
				[8+2*23+2:2*23+2] RoundEP
				[2*23+1:23+1] RoundM
				[23:0] RoundMP
			*/
			pipe_3 = {pipe_2[8 + 23 + 7:8 + 23 + 1], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]} ;
			/* PIPE 4
				[16+4:5] Z
				[4:0] Flags
			*/				
			pipe_4 = {Z_int[32-1:0], Flags_int[4:0]} ;
		end
	end
		
endmodule



module FPMult_PrepModule_dspchain (
		clk,
		rst,
		a,
		b,
		Sa,
		Sb,
		Ea,
		Eb,
		Mp,
		InputExc
	);
	
	// Input ports
	input clk ;
	input rst ;
	input [16-1:0] a ;								// Input A, a 32-bit floating point number
	input [16-1:0] b ;								// Input B, a 32-bit floating point number
	
	// Output ports
	output Sa ;										// A's sign
	output Sb ;										// B's sign
	output [5-1:0] Ea ;								// A's 5
	output [5-1:0] Eb ;								// B's 5
	output [2*10+1:0] Mp ;							// 10 product
	output [4:0] InputExc ;						// Input numbers are exceptions
	
	// Internal signals							// If signal is high...
	wire ANaN ;										// A is a signalling NaN
	wire BNaN ;										// B is a signalling NaN
	wire AInf ;										// A is infinity
	wire BInf ;										// B is infinity
    wire [10-1:0] Ma;
    wire [10-1:0] Mb;
	
	assign ANaN = &(a[16-2:10]) &  |(a[16-2:10]) ;			// All one 5 and not all zero 10 - NaN
	assign BNaN = &(b[16-2:10]) &  |(b[10-1:0]);			// All one 5 and not all zero 10 - NaN
	assign AInf = &(a[16-2:10]) & ~|(a[16-2:10]) ;		// All one 5 and all zero 10 - Infinity
	assign BInf = &(b[16-2:10]) & ~|(b[16-2:10]) ;		// All one 5 and all zero 10 - Infinity
	
	// Check for any exceptions and put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	//assign InputExc = {(ANaN | ANaN | BNaN |BNaN), ANaN, ANaN, BNaN,BNaN} ;
	
	// Take input numbers apart
	assign Sa = a[16-1] ;							// A's sign
	assign Sb = b[16-1] ;							// B's sign
	assign Ea = a[16-2:10];						// Store A's 5 in Ea, unless A is an exception
	assign Eb = b[16-2:10];						// Store B's 5 in Eb, unless B is an exception	
//    assign Ma = a[10_MSB:10_LSB];
  //  assign Mb = b[10_MSB:10_LSB];
	

	// Actual 10 multiplication occurs here
	//assign Mp = ({4'b0001, a[10-1:0]}*{4'b0001, b[10-1:9]}) ;
	assign Mp = ({1'b1,a[10-1:0]}*{1'b1, b[10-1:0]}) ;

	
    //We multiply part of the 10 here
    //Full 10 of A
    //Bits 10_MUL_SPLIT_MSB:10_MUL_SPLIT_LSB of B
   // wire [`ACTUAL_10-1:0] inp_A;
   // wire [`ACTUAL_10-1:0] inp_B;
   // assign inp_A = {1'b1, Ma};
   // assign inp_B = {{(10-(10_MUL_SPLIT_MSB-10_MUL_SPLIT_LSB+1)){1'b0}}, 1'b1, Mb[10_MUL_SPLIT_MSB:10_MUL_SPLIT_LSB]};
   // DW02_mult #(`ACTUAL_10,`ACTUAL_10) u_mult(.A(inp_A), .B(inp_B), .TC(1'b0), .PRODUCT(Mp));
endmodule


module FPMult_ExecuteModule_dspchain(
		a,
		b,
		MpC,
		Ea,
		Eb,
		Sa,
		Sb,
		Sp,
		NormE,
		NormM,
		GRS
    );

	// Input ports
	input [10-1:0] a ;
	input [2*5:0] b ;
	input [2*10+1:0] MpC ;
	input [5-1:0] Ea ;						// A's 5
	input [5-1:0] Eb ;						// B's 5
	input Sa ;								// A's sign
	input Sb ;								// B's sign
	
	// Output ports
	output Sp ;								// Product sign
	output [8:0] NormE ;													// Normalized 5
	output [23-1:0] NormM ;												// Normalized 10
	output GRS ;
	
	wire [2*10+1:0] Mp ;
	
	assign Sp = (Sa ^ Sb) ;												// Equal signs give a positive product
	
   // wire [`ACTUAL_10-1:0] inp_a;
   // wire [`ACTUAL_10-1:0] inp_b;
   // assign inp_a = {1'b1, a};
   // assign inp_b = {{(10-10_MUL_SPLIT_LSB){1'b0}}, 1'b0, b};
   // DW02_mult #(`ACTUAL_10,`ACTUAL_10) u_mult(.A(inp_a), .B(inp_b), .TC(1'b0), .PRODUCT(Mp_temp));
   // DW01_add #(2*`ACTUAL_10) u_add(.A(Mp_temp), .B(MpC<<10_MUL_SPLIT_LSB), .CI(1'b0), .SUM(Mp), .CO());

	//assign Mp = (MpC<<(2*5+1)) + ({4'b0001, a[10-1:0]}*{1'b0, b[2*5:0]}) ;
	assign Mp = MpC;


	assign NormM = (Mp[2*10+1] ? Mp[2*10:0] : Mp[2*10-1:0]); 	// Check for overflow
	assign NormE = (Ea + Eb + Mp[2*10+1]);								// If so, increment 5
	
	assign GRS = ((Mp[10]&(Mp[10+1]))|(|Mp[10-1:0])) ;
	
endmodule

module FPMult_NormalizeModule_dspchain(
		NormM,
		NormE,
		RoundE,
		RoundEP,
		RoundM,
		RoundMP
    );

	// Input Ports
	input [23-1:0] NormM ;									// Normalized 10
	input [8:0] NormE ;									// Normalized 5

	// Output Ports
	output [8:0] RoundE ;
	output [8:0] RoundEP ;
	output [23:0] RoundM ;
	output [23:0] RoundMP ; 
	
// 5 = 5 
// 5 -1 = 4
// NEED to subtract 2^4 -1 = 15

wire [8-1 : 0] bias;

assign bias =  ((1<< (8 -1)) -1);

	assign RoundE = NormE - 9'd15 - 9'd15 + 9'd127 ;
	assign RoundEP = NormE - 9'd15 - 9'd15 + 9'd127 ;
	assign RoundM = NormM ;
	assign RoundMP = NormM ;

endmodule

module FPMult_RoundModule_dspchain(
		RoundM,
		RoundMP,
		RoundE,
		RoundEP,
		Sp,
		GRS,
		InputExc,
		Z,
		Flags
    );

	// Input Ports
	input [23:0] RoundM ;									// Normalized 10
	input [23:0] RoundMP ;									// Normalized 5
	input [8:0] RoundE ;									// Normalized 10 + 1
	input [8:0] RoundEP ;									// Normalized 5 + 1
	input Sp ;												// Product sign
	input GRS ;
	input [4:0] InputExc ;
	
	// Output Ports
	output [32-1:0] Z ;										// Final product
	output [4:0] Flags ;
	
	// Internal Signals
	wire [8:0] FinalE ;									// Rounded 5
	wire [23:0] FinalM;
	wire [23:0] PreShiftM;
	
	assign PreShiftM = GRS ? RoundMP : RoundM ;	// Round up if R and (G or S)
	
	// Post rounding normalization (potential one bit shift> use shifted 10 if there is overflow)
	assign FinalM = (PreShiftM[23] ? {1'b0, PreShiftM[23:1]} : PreShiftM[23:0]) ;
	assign FinalE = (PreShiftM[23] ? RoundEP : RoundE) ; // Increment 5 if a shift was done
	
	
	assign Z = {Sp, FinalE[8-1:0], FinalM[21-1:0], 2'b0} ;   // Putting the pieces together
	assign Flags = InputExc[4:0];

endmodule


module FPAddSub_single_dspchain(
		clk,
		rst,
		a,
		b,
		operation,
		result,
		flags
	);

// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [31:0] a ;								// Input A, a 32-bit floating point number
	input [31:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [31:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754

	reg [68:0]pipe_1;
	reg [54:0]pipe_2;
	reg [45:0]pipe_3;


//internal module wires

//output ports
	wire Opout;
	wire Sa;
	wire Sb;
	wire MaxAB;
	wire [7:0] CExp;
	wire [4:0] Shift;
	wire [22:0] Mmax;
	wire [4:0] InputExc;
	wire [23:0] Mmin_3;

	wire [32:0] SumS_5 ;
	wire [4:0] Shift_1;							
	wire PSgn ;							
	wire Opr ;	
	
	wire [22:0] NormM ;				// Normalized mantissa
	wire [8:0] NormE ;					// Adjusted exponent
	wire ZeroSum ;						// Zero flag
	wire NegE ;							// Flag indicating negative exponent
	wire R ;								// Round bit
	wire S ;								// Final sticky bit
	wire FG ;

FPAddSub_a_dspchain M1(a,b,operation,Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3);

FpAddSub_b_dspchain M2(pipe_1[51:29],pipe_1[23:0],pipe_1[67],pipe_1[66],pipe_1[65],pipe_1[68],SumS_5,Shift_1,PSgn,Opr);

FPAddSub_c_dspchain M3(pipe_2[54:22],pipe_2[21:17],pipe_2[16:9],NormM,NormE,ZeroSum,NegE,R,S,FG);

FPAddSub_d_dspchain M4(pipe_3[13],pipe_3[22:14],pipe_3[45:23],pipe_3[11],pipe_3[10],pipe_3[9],pipe_3[8],pipe_3[7],pipe_3[6],pipe_3[5],pipe_3[12],pipe_3[4:0],result,flags );


always @ (posedge clk) begin	
		if(rst) begin
			pipe_1 <= 0;
			pipe_2 <= 0;
			pipe_3 <= 0;
		end 
		else begin
/*
pipe_1:
	[68] Opout;
	[67] Sa;
	[66] Sb;
	[65] MaxAB;
	[64:57] CExp;
	[56:52] Shift;
	[51:29] Mmax;
	[28:24] InputExc;
	[23:0] Mmin_3;	
*/

pipe_1 <= {Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3};

/*
pipe_2:
	[54:22]SumS_5;
	[21:17]Shift;
	[16:9]CExp;	
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_2 <= {SumS_5,Shift_1,pipe_1[64:57], pipe_1[67], pipe_1[66], pipe_1[68], pipe_1[65], pipe_1[28:24] };

/*
pipe_3:
	[45:23] NormM ;				
	[22:14] NormE ;					
	[13]ZeroSum ;						
	[12]NegE ;							
	[11]R ;								
	[10]S ;								
	[9]FG ;
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_3 <= {NormM,NormE,ZeroSum,NegE,R,S,FG, pipe_2[8], pipe_2[7], pipe_2[6], pipe_2[5], pipe_2[4:0] };

end
end

endmodule

// Prealign + Align + Shift 1 + Shift 2
module FPAddSub_a_dspchain(
		A,
		B,
		operation,
		Opout,
		Sa,
		Sb,
		MaxAB,
		CExp,
		Shift,
		Mmax,
		InputExc,
		Mmin_3
		
		
	);
	
	// Input ports
	input [31:0] A ;										// Input A, a 32-bit floating point number
	input [31:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	//output ports
	output Opout;
	output Sa;
	output Sb;
	output MaxAB;
	output [7:0] CExp;
	output [4:0] Shift;
	output [22:0] Mmax;
	output [4:0] InputExc;
	output [23:0] Mmin_3;	
							
	wire [9:0] ShiftDet ;							
	wire [30:0] Aout ;
	wire [30:0] Bout ;
	

	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [7:0] DAB ;										// ExpA - ExpB					
	wire [7:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[30:23]) & |(A[22:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[30:23]) & |(B[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[30:23]) & ~|(A[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[30:23]) & ~|(B[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
  assign DAB = (A[30:23] + ~(B[30:23]) + 1) ;
	assign DBA = (B[30:23] + ~(A[30:23]) + 1) ;

	assign Sa = A[31] ;									// A's sign bit
	assign Sb = B[31] ;									// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[30:0] ;
	assign Bout = B[30:0] ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Output ports
													// Number of steps to smaller mantissa shift right
	wire [22:0] Mmin_1 ;							// Smaller mantissa 
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (Aout[30:0] < Bout[30:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[9:5] : ShiftDet[4:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin_1 = MaxAB ? Aout[22:0] : Bout[22:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? Bout[22:0]: Aout[22:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? Bout[30:23] : Aout[30:23]) ;	

// Input ports
					// Smaller mantissa after 16|12|8|4 shift
	wire [2:0] Shift_1 ;						// Shift amount
	
	assign Shift_1 = Shift [4:2];

	wire [23:0] Mmin_2 ;						// The smaller mantissa
	
	// Internal signals
	reg	  [23:0]		Lvl1;
	reg	  [23:0]		Lvl2;
	wire    [47:0]    Stage1;	
	integer           i;                // Loop variable
	
	always @(*) begin						
		// Rotate by 16?
		Lvl1 <= Shift_1[2] ? {17'b00000000000000001, Mmin_1[22:16]} : {1'b1, Mmin_1}; 
	end
	
	assign Stage1 = {Lvl1, Lvl1};
	
	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift_1[1:0])
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[23:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[23:19] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[23:15] <= 0; end
			// Rotate by 12	
			2'b11:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[23:11] <= 0; end
	  endcase
	end
	
	// Assign output to next shift stage
	assign Mmin_2 = Lvl2;
								// Smaller mantissa after 16|12|8|4 shift
	wire [1:0] Shift_2 ;						// Shift amount
	
	assign Shift_2 =Shift  [1:0] ;
					// The smaller mantissa
	
	// Internal Signal
	reg	  [23:0]		Lvl3;
	wire    [47:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {Mmin_2, Mmin_2};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_2[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[23:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[23] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[23:22] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[23:21] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin_3 = Lvl3;	

	
endmodule

module FpAddSub_b_dspchain(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		SumS_5,
		Shift,
		PSgn,
		Opr
);
	input [22:0] Mmax ;					// The larger mantissa
	input [23:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	wire [32:0] Sum ;	
						// Output ports
	output [32:0] SumS_5 ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount				// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation

	// Perform effective operation
	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, 8'b00000000} - {Mmin, 8'b00000000}) : ({1'b1, Mmax, 8'b00000000} + {Mmin, 8'b00000000}) ;
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

		// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[32] ? 5'b00000 :	 
		Sum[31] ? 5'b00001 : 
		Sum[30] ? 5'b00010 : 
		Sum[29] ? 5'b00011 : 
		Sum[28] ? 5'b00100 : 
		Sum[27] ? 5'b00101 : 
		Sum[26] ? 5'b00110 : 
		Sum[25] ? 5'b00111 :
		Sum[24] ? 5'b01000 :
		Sum[23] ? 5'b01001 :
		Sum[22] ? 5'b01010 :
		Sum[21] ? 5'b01011 :
		Sum[20] ? 5'b01100 :
		Sum[19] ? 5'b01101 :
		Sum[18] ? 5'b01110 :
		Sum[17] ? 5'b01111 :
		Sum[16] ? 5'b10000 :
		Sum[15] ? 5'b10001 :
		Sum[14] ? 5'b10010 :
		Sum[13] ? 5'b10011 :
		Sum[12] ? 5'b10100 :
		Sum[11] ? 5'b10101 :
		Sum[10] ? 5'b10110 :
		Sum[9] ? 5'b10111 :
		Sum[8] ? 5'b11000 :
		Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [32:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[16:0], 16'b0000000000000000} : Sum; 
	end
	
	// Assign outputs
	assign SumS_5 = Lvl1;	

endmodule

module FPAddSub_c_dspchain(
		SumS_5,
		Shift,
		CExp,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [32:0] SumS_5 ;						// Smaller mantissa after 16|12|8|4 shift
	
	input [4:0] Shift ;						// Shift amount
	
// Input ports
	
	input [7:0] CExp ;
	

	// Output ports
	output [22:0] NormM ;				// Normalized mantissa
	output [8:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;


	wire [3:0]Shift_1;
	assign Shift_1 = Shift [3:0];
	// Output ports
	wire [32:0] SumS_7 ;						// The smaller mantissa
	
	reg	  [32:0]		Lvl2;
	wire    [65:0]    Stage1;	
	reg	  [32:0]		Lvl3;
	wire    [65:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {SumS_5, SumS_5};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[32:0];       		
			// Rotate by 4
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_1[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[32:0];
			// Rotate by 1
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign SumS_7 = Lvl3;						// Take out smaller mantissa



	
	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [8:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [8:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = SumS_7[32] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|SumS_7 ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[8] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = SumS_7[31:9] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = SumS_7[8] ; 
	assign R = SumS_7[7] ;
	assign S = |SumS_7[6:0] ;		
	
endmodule

module FPAddSub_d_dspchain(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		NegE,
		InputExc,
		P,
		Flags 
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [8:0] NormE ;				// Normalized exponent
	input [22:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	

	input NegE ;						// Negative exponent?
	input [4:0] InputExc ;					// Exceptions in inputs A and B

	// Output ports
	output [31:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// 
	wire [31:0] Z ;					// Final result
	wire EOF ;
	
	// Internal signals
	wire [23:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [22:0] RoundM ;				// The final rounded sum
	wire [8:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	wire FSgn;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[22:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[23] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? 8'b00000000 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[7:0], RoundM[22:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[8];

/////////////////////////////////////////////////////////////////////////////////////////////////////////



	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[30:23]) & ~|(Z[30:23]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule

`endif 


module spram_2048_40bit (
    clk,
    address,
    wren,
    data,
    out
);
parameter AWIDTH=11;
parameter NUM_WORDS=2048;
parameter DWIDTH=40;
input clk;
input [(AWIDTH-1):0] address;
input  wren;
input [(DWIDTH-1):0] data;
output reg [(DWIDTH-1):0] out;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren) begin
      ram[address] <= data;
  end
  else begin
      out <= ram[address];
  end
end
  
`else

defparam u_single_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_single_port_ram.DATA_WIDTH = DWIDTH;

single_port_ram u_single_port_ram(
.addr(address),
.we(wren),
.data(data),
.out(out),
.clk(clk)
);

`endif

endmodule

`timescale 1ns / 1ps


`define BFLOAT16
`ifdef BFLOAT16
`define EXPONENT 8
`define MANTISSA 7
`else // for ieee half precision fp16
`define EXPONENT 5
`define MANTISSA 10
`endif

`define SIGN 1
`define DWIDTH (`SIGN+`EXPONENT+`MANTISSA)

module tensor_block_bf16(
	clk,
	reset,
	
	data_in,
	cascade_in,
	acc0_in,
	acc1_in,
	acc2_in,
	accumulator_input1_select,

	out0,
	out1,
	out2,
	cascade_out,
	acc0_out,
	acc1_out,
	acc2_out,

	mux1_select,
	dot_unit_input_1_enable,
	bank0_data_in_enable,
	bank1_data_in_enable,
	cascade_out_select,
	dot_unit_input_2_select

	);

input 	[79:0] data_in;
input	[79:0] cascade_in;
input	[31:0] acc0_in;
input	[31:0] acc1_in;
input	[31:0] acc2_in;
input 	[2:0] accumulator_input1_select;


output	[31:0] out0;
output	[31:0] out1;
output	[31:0] out2;
output	[79:0] cascade_out;
output	[31:0] acc0_out;
output	[31:0] acc1_out;
output	[31:0] acc2_out;

//Inputs to take into account
input clk;
input reset;

// Logic to be created for 
input mux1_select;
input dot_unit_input_1_enable;
input bank0_data_in_enable;
input bank1_data_in_enable;
input cascade_out_select;
input dot_unit_input_2_select;


wire [79:0]mux1_out;
assign mux1_out = mux1_select ? cascade_in : data_in;

reg [79:0]dot_unit_input_1;

// D Flip Flop with reset and enable
always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) dot_unit_input_1 <= 0;
	else if (dot_unit_input_1_enable) dot_unit_input_1 <= data_in;
end

// Register Bank 0 
reg[79:0] bank0_reg0;
reg[79:0] bank0_reg1;
reg[79:0] bank0_reg2;

always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) begin
		bank0_reg0 <= 0;
		bank0_reg1 <= 0;
		bank0_reg2 <= 0;
	end
	else if (bank0_data_in_enable) begin
		bank0_reg0 <= mux1_out;
		bank0_reg1 <= bank0_reg0;
		bank0_reg2 <= bank0_reg1;
	end
end

// Register Bank 1 
reg[79:0] bank1_reg0;
reg[79:0] bank1_reg1;
reg[79:0] bank1_reg2;

always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) begin
		bank1_reg0 <= 0;
		bank1_reg1 <= 0;
		bank1_reg2 <= 0;
	end
	else if (bank1_data_in_enable) begin
		bank1_reg0 <= mux1_out;
		bank1_reg1 <= bank0_reg0;
		bank1_reg2 <= bank0_reg1;
	end
end

// Output cascade out
assign cascade_out = cascade_out_select ? bank1_reg2 : bank0_reg2;

// Providing second input to all 3 dot product units
wire [79:0]dot_unit_input_2_0;
wire [79:0]dot_unit_input_2_1;
wire [79:0]dot_unit_input_2_2;

assign dot_unit_input_2_0 = dot_unit_input_2_select ? bank1_reg0 : bank0_reg0;
assign dot_unit_input_2_1 = dot_unit_input_2_select ? bank1_reg1 : bank0_reg1;
assign dot_unit_input_2_2 = dot_unit_input_2_select ? bank1_reg2 : bank0_reg2;

wire [31:0] dot_unit_output_0;
wire [31:0] dot_unit_output_1;
wire [31:0] dot_unit_output_2;

dot_product_unit dot_unit0 (clk, reset, dot_unit_input_1, dot_unit_input_2_0, dot_unit_output_0);
dot_product_unit dot_unit1 (clk, reset, dot_unit_input_1, dot_unit_input_2_1, dot_unit_output_1);
dot_product_unit dot_unit2 (clk, reset, dot_unit_input_1, dot_unit_input_2_2, dot_unit_output_2);

// Flopping after dot product compute
reg [31:0] dot_unit_output_0_flopped;
reg [31:0] dot_unit_output_1_flopped;
reg [31:0] dot_unit_output_2_flopped;

always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) begin
		dot_unit_output_0_flopped <= 0;
		dot_unit_output_1_flopped <= 0;
		dot_unit_output_2_flopped <= 0;
	end
	else begin
		dot_unit_output_0_flopped <= dot_unit_output_0;
		dot_unit_output_1_flopped <= dot_unit_output_1;
		dot_unit_output_2_flopped <= dot_unit_output_2;
	end
end

wire [31:0] accumulator_unit0_input1;
wire [31:0] accumulator_unit1_input1;
wire [31:0] accumulator_unit2_input1;

wire [31:0] accumulator_unit_output_0;
wire [31:0] accumulator_unit_output_1;
wire [31:0] accumulator_unit_output_2;

reg [31:0] accumulator_unit_output_0_flopped;
reg [31:0] accumulator_unit_output_1_flopped;
reg [31:0] accumulator_unit_output_2_flopped;

reg [31:0] acc0_in_flopped;
reg [31:0] acc1_in_flopped;
reg [31:0] acc2_in_flopped;

// 3 mux's for selecting acc_in or acc_out_flopped
assign accumulator_unit0_input1 = accumulator_input1_select[0] ?  accumulator_unit_output_0_flopped : acc0_in_flopped;
assign accumulator_unit1_input1 = accumulator_input1_select[1] ?  accumulator_unit_output_1_flopped : acc1_in_flopped;
assign accumulator_unit2_input1 = accumulator_input1_select[2] ?  accumulator_unit_output_2_flopped : acc2_in_flopped;

// Flopping the accumulator outputs and acc_in 
always @ (posedge clk, posedge reset) begin
	if (reset == 1'b1) begin
		accumulator_unit_output_0_flopped <= 0;
		accumulator_unit_output_1_flopped <= 0;
		accumulator_unit_output_2_flopped <= 0;
		acc0_in_flopped <= 0;
		acc1_in_flopped <= 0;
		acc2_in_flopped <= 0;
	end
	else begin
		accumulator_unit_output_0_flopped <= accumulator_unit_output_0;
		accumulator_unit_output_1_flopped <= accumulator_unit_output_1;
		accumulator_unit_output_2_flopped <= accumulator_unit_output_2;
		acc0_in_flopped <= acc0_in;
		acc1_in_flopped <= acc1_in;
		acc2_in_flopped <= acc2_in;
	end
end

// Accumulator units
accumulator acc_unit0 (clk, reset, dot_unit_output_0_flopped, accumulator_unit0_input1, accumulator_unit_output_0 );
accumulator acc_unit1 (clk, reset, dot_unit_output_1_flopped, accumulator_unit1_input1, accumulator_unit_output_1 );
accumulator acc_unit2 (clk, reset, dot_unit_output_2_flopped, accumulator_unit2_input1, accumulator_unit_output_2 );

assign acc0_out = accumulator_unit_output_0;
assign acc1_out = accumulator_unit_output_1;
assign acc2_out = accumulator_unit_output_2;

//Taking the top 25 bits from the 32 bit accumulation number
assign out0= accumulator_unit_output_0;
assign out1= accumulator_unit_output_1;
assign out2= accumulator_unit_output_2;

endmodule

module dot_product_unit (
	clk,
	reset,
	data_in_1,
	data_in_2,
	data_out
	);
input clk;
input reset;
input [79:0] data_in_1;
input [79:0] data_in_2;
output [31:0] data_out;

wire [15:0] mult1_in1;
wire [15:0] mult1_in2;
wire [31:0] mult1_out;
wire [15:0] mult2_in1;
wire [15:0] mult2_in2;
wire [31:0] mult2_out;
wire [15:0] mult3_in1;
wire [15:0] mult3_in2;
wire [31:0] mult3_out;
wire [15:0] mult4_in1;
wire [15:0] mult4_in2;
wire [31:0] mult4_out;
wire [15:0] mult5_in1;
wire [15:0] mult5_in2;
wire [31:0] mult5_out;
reg [31:0] mult1_out_reg;
reg [31:0] mult2_out_reg;
reg [31:0] mult3_out_reg;
reg [31:0] mult4_out_reg;
reg [31:0] mult5_out_reg;

wire [4:0] flags_dummy_1;
wire [4:0] flags_dummy_2;
wire [4:0] flags_dummy_3;
wire [4:0] flags_dummy_4;
wire [4:0] flags_dummy_5;

assign mult1_in1 = data_in_1[15:0];
assign mult1_in2 = data_in_2[15:0];
FPMult_16 mult_1_dut(clk,reset,mult1_in1,mult1_in2,mult1_out,flags_dummy_1);


assign mult2_in1 = data_in_1[31:16];
assign mult2_in2 = data_in_2[31:16];
FPMult_16 mult_2_dut(clk,reset,mult2_in1,mult2_in2,mult2_out,flags_dummy_2);

assign mult3_in1 = data_in_1[47:32];
assign mult3_in2 = data_in_2[47:32];
FPMult_16 mult_3_dut(clk,reset,mult3_in1,mult3_in2,mult3_out,flags_dummy_3);

assign mult4_in1 = data_in_1[63:48];
assign mult4_in2 = data_in_2[63:48];
FPMult_16 mult_4_dut(clk,reset,mult4_in1,mult4_in2,mult4_out,flags_dummy_4);

assign mult5_in1 = data_in_1[79:54];
assign mult5_in2 = data_in_2[79:54];
FPMult_16 mult_5_dut(clk,reset,mult5_in1,mult5_in2,mult5_out,flags_dummy_5);

always@(posedge clk) begin 
mult1_out_reg <= mult1_out; 
mult2_out_reg <= mult2_out; 
mult3_out_reg <= mult3_out; 
mult4_out_reg <= mult4_out; 
mult5_out_reg <= mult5_out; 
end

sum_5_times sum_it_up(clk, reset, mult1_out_reg, mult2_out_reg, mult3_out_reg, mult4_out_reg, mult5_out_reg, data_out);
//assign data_out = 	mult1_out + mult2_out + mult3_out + mult4_out + mult5_out +  
//					mult6_out + mult7_out + mult8_out + mult9_out + mult10_out;
endmodule


module sum_5_times (clk, reset, num1, num2, num3, num4, num5, out);

input clk;
input reset;
input [31:0]num1;
input [31:0]num2;
input [31:0]num3;
input [31:0]num4;
input [31:0]num5;
output [31:0] out;

wire [31:0]add_1_out;
wire [31:0]add_2_out;
wire [31:0]add_3_out;
wire [31:0]add_4_out;

reg [31:0] add_1_out_reg; 
reg [31:0] add_2_out_reg;
reg [31:0] add_3_out_reg;

wire [4:0] dummy_flag_1;
wire [4:0] dummy_flag_2;
wire [4:0] dummy_flag_3;
wire [4:0] dummy_flag_4;


FPAddSub_single_32 sum_10_times_adder_1(clk,reset,num1,num2,1'b0,add_1_out,dummy_flag_1);
always@(posedge clk) begin 
add_1_out_reg<= add_1_out;
end

FPAddSub_single_32 sum_10_times_adder_2(clk,reset,num3,num4,1'b0,add_2_out,dummy_flag_2);
always@(posedge clk) begin 
add_2_out_reg<= add_2_out;
end

FPAddSub_single_32 sum_10_times_adder_3(clk,reset,add_1_out_reg,add_2_out_reg,1'b0,add_3_out,dummy_flag_3);
always@(posedge clk) begin 
add_3_out_reg<= add_3_out;
end
reg [31:0] num5_del0,num5_del1;

always@(posedge clk) begin 
num5_del0<= num5;
num5_del1<= num5_del0;
end

FPAddSub_single_32 sum_10_times_adder_4(clk,reset,add_3_out_reg,num5_del1,1'b0,add_4_out,dummy_flag_4);

assign out = add_4_out;

endmodule

module accumulator (
	clk,
	reset,
	input_accumlator_1,
	input_accumlator_2,
	output_accumlator
	);
input clk;
input reset;
input [31:0] input_accumlator_1;
input [31:0] input_accumlator_2;
output [31:0] output_accumlator;

wire [4:0] flags; //dummy

FPAddSub_single_32 accumulator_definition(
		clk,
		reset,
		input_accumlator_1,
		input_accumlator_2,
		1'b0,			// 0 add, 1 sub
		output_accumlator,
		flags
	);

endmodule


module FPAddSub_single_32(
		clk,
		rst,
		a,
		b,
		operation,
		result,
		flags
	);

  // Clock and reset
  	input clk ;										// Clock signal
  	input rst ;										// Reset (active high, resets pipeline registers)
  	
  	// Input ports
  	input [31:0] a ;								// Input A, a 32-bit floating point number
  	input [31:0] b ;								// Input B, a 32-bit floating point number
  	input operation ;								// Operation select signal
  	
  	// Output ports
  	output [31:0] result ;						// Result of the operation
  	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754
  
  	reg [68:0]pipe_1;
  	reg [54:0]pipe_2;
  	reg [45:0]pipe_3;
  
  
  //internal module wires
  
  //output ports
  	wire Opout;
  	wire Sa;
  	wire Sb;
  	wire MaxAB;
  	wire [7:0] CExp;
  	wire [4:0] Shift;
  	wire [22:0] Mmax;
  	wire [4:0] InputExc;
  	wire [23:0] Mmin_3;
  
  	wire [32:0] SumS_5 ;
  	wire [4:0] Shift_1;							
  	wire PSgn ;							
  	wire Opr ;	
  	
  	wire [22:0] NormM ;				// Normalized mantissa
  	wire [8:0] NormE ;					// Adjusted exponent
  	wire ZeroSum ;						// Zero flag
  	wire NegE ;							// Flag indicating negative exponent
  	wire R ;								// Round bit
  	wire S ;								// Final sticky bit
  	wire FG ;
  
  FPAddSub_a_32 M1(a,b,operation,Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3);
  
  FpAddSub_b_32 M2(pipe_1[51:29],pipe_1[23:0],pipe_1[67],pipe_1[66],pipe_1[65],pipe_1[68],SumS_5,Shift_1,PSgn,Opr);
  
  FPAddSub_c_32 M3(pipe_2[54:22],pipe_2[21:17],pipe_2[16:9],NormM,NormE,ZeroSum,NegE,R,S,FG);
  
  FPAddSub_d_32 M4(pipe_3[13],pipe_3[22:14],pipe_3[45:23],pipe_3[11],pipe_3[10],pipe_3[9],pipe_3[8],pipe_3[7],pipe_3[6],pipe_3[5],pipe_3[12],pipe_3[4:0],result,flags );
  
  
  always @ (posedge clk) begin	
  		if(rst) begin
  			pipe_1 <= 0;
  			pipe_2 <= 0;
  			pipe_3 <= 0;
  		end 
  		else begin
  /*
  pipe_1:
  	[68] Opout;
  	[67] Sa;
  	[66] Sb;
  	[65] MaxAB;
  	[64:57] CExp;
  	[56:52] Shift;
  	[51:29] Mmax;
  	[28:24] InputExc;
  	[23:0] Mmin_3;	
  */
  
  pipe_1 <= {Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3};
  
  /*
  pipe_2:
  	[54:22]SumS_5;
  	[21:17]Shift;
  	[16:9]CExp;	
  	[8]Sa;
  	[7]Sb;
  	[6]operation;
  	[5]MaxAB;	
  	[4:0]InputExc
  */
  
  pipe_2 <= {SumS_5,Shift_1,pipe_1[64:57], pipe_1[67], pipe_1[66], pipe_1[68], pipe_1[65], pipe_1[28:24] };
  
  /*
  pipe_3:
  	[45:23] NormM ;				
  	[22:14] NormE ;					
  	[13]ZeroSum ;						
  	[12]NegE ;							
  	[11]R ;								
  	[10]S ;								
  	[9]FG ;
  	[8]Sa;
  	[7]Sb;
  	[6]operation;
  	[5]MaxAB;	
  	[4:0]InputExc
  */
  
  pipe_3 <= {NormM,NormE,ZeroSum,NegE,R,S,FG, pipe_2[8], pipe_2[7], pipe_2[6], pipe_2[5], pipe_2[4:0] };
  
  end
  end


endmodule

module FPAddSub_a_32(
		A,
		B,
		operation,
		Opout,
		Sa,
		Sb,
		MaxAB,
		CExp,
		Shift,
		Mmax,
		InputExc,
		Mmin_3
		
		
	);
	
	// Input ports
	input [31:0] A ;										// Input A, a 32-bit floating point number
	input [31:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	//output ports
	output Opout;
	output Sa;
	output Sb;
	output MaxAB;
	output [7:0] CExp;
	output [4:0] Shift;
	output [22:0] Mmax;
	output [4:0] InputExc;
	output [23:0] Mmin_3;	
							
	wire [9:0] ShiftDet ;							
	wire [30:0] Aout ;
	wire [30:0] Bout ;
	

	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [7:0] DAB ;										// ExpA - ExpB					
	wire [7:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[30:23]) & |(A[22:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[30:23]) & |(B[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[30:23]) & ~|(A[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[30:23]) & ~|(B[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
	assign DAB = (A[30:23] + ~(B[30:23]) + 1) ;
	assign DBA = (B[30:23] + ~(A[30:23]) + 1) ;
	
	assign Sa = A[31] ;									// A's sign bit
	assign Sb = B[31] ;									// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[30:0] ;
	assign Bout = B[30:0] ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Output ports
													// Number of steps to smaller mantissa shift right
	wire [22:0] Mmin_1 ;							// Smaller mantissa 
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (Aout[30:0] < Bout[30:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[9:5] : ShiftDet[4:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin_1 = MaxAB ? Aout[22:0] : Bout[22:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? Bout[22:0]: Aout[22:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? Bout[30:23] : Aout[30:23]) ;	

// Input ports
					// Smaller mantissa after 16|12|8|4 shift
	wire [2:0] Shift_1 ;						// Shift amount
	
	assign Shift_1 = Shift [4:2];

	wire [23:0] Mmin_2 ;						// The smaller mantissa
	
	// Internal signals
	reg	  [23:0]		Lvl1;
	reg	  [23:0]		Lvl2;
	wire    [47:0]    Stage1;	
	integer           i;                // Loop variable
	
	always @(*) begin						
		// Rotate by 16?
		Lvl1 <= Shift_1[2] ? {17'b00000000000000001, Mmin_1[22:16]} : {1'b1, Mmin_1}; 
	end
	
	assign Stage1 = {Lvl1, Lvl1};
	
	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift_1[1:0])
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[23:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[23:19] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[23:15] <= 0; end
			// Rotate by 12	
			2'b11:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[23:11] <= 0; end
	  endcase
	end
	
	// Assign output to next shift stage
	assign Mmin_2 = Lvl2;
								// Smaller mantissa after 16|12|8|4 shift
	wire [1:0] Shift_2 ;						// Shift amount
	
	assign Shift_2 =Shift  [1:0] ;
					// The smaller mantissa
	
	// Internal Signal
	reg	  [23:0]		Lvl3;
	wire    [47:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {Mmin_2, Mmin_2};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_2[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[23:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[23] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[23:22] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[23:21] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin_3 = Lvl3;	

	
endmodule

module FpAddSub_b_32(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		SumS_5,
		Shift,
		PSgn,
		Opr
);
	input [22:0] Mmax ;					// The larger mantissa
	input [23:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	wire [32:0] Sum ;	
						// Output ports
	output [32:0] SumS_5 ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount				// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation

	// Perform effective operation
	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, 8'b00000000} - {Mmin, 8'b00000000}) : ({1'b1, Mmax, 8'b00000000} + {Mmin, 8'b00000000}) ;
	
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

		// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[32] ? 5'b00000 :	 
		Sum[31] ? 5'b00001 : 
		Sum[30] ? 5'b00010 : 
		Sum[29] ? 5'b00011 : 
		Sum[28] ? 5'b00100 : 
		Sum[27] ? 5'b00101 : 
		Sum[26] ? 5'b00110 : 
		Sum[25] ? 5'b00111 :
		Sum[24] ? 5'b01000 :
		Sum[23] ? 5'b01001 :
		Sum[22] ? 5'b01010 :
		Sum[21] ? 5'b01011 :
		Sum[20] ? 5'b01100 :
		Sum[19] ? 5'b01101 :
		Sum[18] ? 5'b01110 :
		Sum[17] ? 5'b01111 :
		Sum[16] ? 5'b10000 :
		Sum[15] ? 5'b10001 :
		Sum[14] ? 5'b10010 :
		Sum[13] ? 5'b10011 :
		Sum[12] ? 5'b10100 :
		Sum[11] ? 5'b10101 :
		Sum[10] ? 5'b10110 :
		Sum[9] ? 5'b10111 :
		Sum[8] ? 5'b11000 :
		Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [32:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[16:0], 16'b0000000000000000} : Sum; 
	end
	
	// Assign outputs
	assign SumS_5 = Lvl1;	

endmodule

module FPAddSub_c_32(
		SumS_5,
		Shift,
		CExp,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [32:0] SumS_5 ;						// Smaller mantissa after 16|12|8|4 shift
	
	input [4:0] Shift ;						// Shift amount
	
// Input ports
	
	input [7:0] CExp ;
	

	// Output ports
	output [22:0] NormM ;				// Normalized mantissa
	output [8:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;


	wire [3:0]Shift_1;
	assign Shift_1 = Shift [3:0];
	// Output ports
	wire [32:0] SumS_7 ;						// The smaller mantissa
	
	reg	  [32:0]		Lvl2;
	wire    [65:0]    Stage1;	
	reg	  [32:0]		Lvl3;
	wire    [65:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {SumS_5, SumS_5};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[32:0];       		
			// Rotate by 4
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_1[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[32:0];
			// Rotate by 1
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign SumS_7 = Lvl3;						// Take out smaller mantissa



	
	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [8:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [8:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = SumS_7[32] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|SumS_7 ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[8] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	


	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = SumS_7[31:9] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = SumS_7[8] ; 
	assign R = SumS_7[7] ;
	assign S = |SumS_7[6:0] ;		
	
endmodule

module FPAddSub_d_32(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		NegE,
		InputExc,
		P,
		Flags 
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [8:0] NormE ;				// Normalized exponent
	input [22:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	

	input NegE ;						// Negative exponent?
	input [4:0] InputExc ;					// Exceptions in inputs A and B

	// Output ports
	output [31:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// 
	wire [31:0] Z ;					// Final result
	wire EOF ;
	
	// Internal signals
	wire [23:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [22:0] RoundM ;				// The final rounded sum
	wire [8:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	wire FSgn;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[22:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[23] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? 8'b00000000 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[7:0], RoundM[22:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[8];

/////////////////////////////////////////////////////////////////////////////////////////////////////////



	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[30:23]) & ~|(Z[30:23]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule

//////////////////////////////////////////////////////////////////////////////////
//
// Module Name:    FPMult
//
//////////////////////////////////////////////////////////////////////////////////

module FPMult_16(
		clk,
		rst,
		a,
		b,
		result,
		flags
    );
	
	// Input Ports
	input clk ;							// Clock
	input rst ;							// Reset signal
	input [16-1:0] a;						// Input A, a 32-bit floating point number
	input [16-1:0] b;						// Input B, a 32-bit floating point number
	
	// Output ports
	output [32-1:0] result ;					// Product, result of the operation, 32-bit FP number
	output [4:0] flags ;						// Flags indicating exceptions according to IEEE754
	
	// Internal signals
	wire [32-1:0] Z_int ;					// Product, result of the operation, 32-bit FP number
	wire [4:0] Flags_int ;						// Flags indicating exceptions according to IEEE754
	
	wire Sa ;							// A's sign
	wire Sb ;							// B's sign
	wire Sp ;							// Product sign
	wire [8-1:0] Ea ;					// A's exponent
	wire [8-1:0] Eb ;					// B's exponent
	wire [2*7+1:0] Mp ;					// Product 7
	wire [4:0] InputExc ;						// Exceptions in inputs
	wire [23-1:0] NormM ;					// Normalized 7
	wire [8:0] NormE ;					// Normalized exponent
	wire [23:0] RoundM ;					// Normalized 7
	wire [8:0] RoundE ;					// Normalized exponent
	wire [23:0] RoundMP ;					// Normalized 7
	wire [8:0] RoundEP ;					// Normalized exponent
	wire GRS ;

	//reg [63:0] pipe_0;						// Pipeline register Input->Prep
	reg [2*16-1:0] pipe_0;					// Pipeline register Input->Prep

	//reg [92:0] pipe_1;						// Pipeline register Prep->Execute
	//reg [3*7+2*8+7:0] pipe_1;			// Pipeline register Prep->Execute
	reg [3*7+2*8+18:0] pipe_1;

	//reg [38:0] pipe_2;						// Pipeline register Execute->Normalize
	reg [23+8+7:0] pipe_2;				// Pipeline register Execute->Normalize
	
	//reg [72:0] pipe_3;						// Pipeline register Normalize->Round
	reg [2*23+2*8+10:0] pipe_3;			// Pipeline register Normalize->Round

	//reg [36:0] pipe_4;						// Pipeline register Round->Output
	reg [32+4:0] pipe_4;					// Pipeline register Round->Output
	
	assign result = pipe_4[32+4:5] ;
	assign flags = pipe_4[4:0] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPMult_PrepModule PrepModule(clk, rst, pipe_0[2*16-1:16], pipe_0[16-1:0], Sa, Sb, Ea[8-1:0], Eb[8-1:0], Mp[2*7+1:0], InputExc[4:0]) ;

	// Perform (unsigned) 7 multiplication
	FPMult_ExecuteModule ExecuteModule(pipe_1[3*7+8*2+7:2*7+2*8+8], pipe_1[2*7+2*8+7:2*7+7], pipe_1[2*7+6:5], pipe_1[2*7+2*8+6:2*7+8+7], pipe_1[2*7+8+6:2*7+7], pipe_1[2*7+2*8+8], pipe_1[2*7+2*8+7], Sp, NormE[8:0], NormM[23-1:0], GRS) ;

	// Round result and if necessary, perform a second (post-rounding) normalization step
	FPMult_NormalizeModule NormalizeModule(pipe_2[23-1:0], pipe_2[23+8:23], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]) ;		

	// Round result and if necessary, perform a second (post-rounding) normalization step
	//FPMult_RoundModule RoundModule(pipe_3[47:24], pipe_3[23:0], pipe_3[65:57], pipe_3[56:48], pipe_3[66], pipe_3[67], pipe_3[72:68], Z_int[31:0], Flags_int[4:0]) ;		
	FPMult_RoundModule RoundModule(pipe_3[2*23+1:23+1], pipe_3[23:0], pipe_3[2*23+2*8+3:2*23+8+3], pipe_3[2*23+8+2:2*23+2], pipe_3[2*23+2*8+4], pipe_3[2*23+2*8+5], pipe_3[2*23+2*8+10:2*23+2*8+6], Z_int[32-1:0], Flags_int[4:0]) ;		

				
//adding always@ (*) instead of posedge clock to make design combinational
	always @ (*) begin	
		if(rst) begin
			pipe_0 = 0;
			pipe_1 = 0;
			pipe_2 = 0; 
			pipe_3 = 0;
			pipe_4 = 0;
		end 
		else begin		
			/* PIPE 0
				[2*16-1:16] A
				[16-1:0] B
			*/
                       pipe_0 = {a, b} ;


			/* PIPE 1
				[2*8+3*7 + 18: 2*8+2*7 + 18] //pipe_0[16+7-1:16] , 7 of A
				[2*8+2*7 + 17 :2*8+2*7 + 9] // pipe_0[8:0]
				[2*8+2*7 + 8] Sa
				[2*8+2*7 + 7] Sb
				[2*8+2*7 + 6:8+2*7+7] Ea
				[8+2*7+6:2*7+7] Eb
				[2*7+1+5:5] Mp
				[4:0] InputExc
			*/
			//pipe_1 <= {pipe_0[16+7-1:16], pipe_0[7_MUL_SPLIT_LSB-1:0], Sa, Sb, Ea[8-1:0], Eb[8-1:0], Mp[2*7-1:0], InputExc[4:0]} ;
			pipe_1 = {pipe_0[16+7-1:16], pipe_0[8:0], Sa, Sb, Ea[8-1:0], Eb[8-1:0], Mp[2*7+1:0], InputExc[4:0]} ;
			
			/* PIPE 2
				[8+ 23 + 7:8+ 23 + 3] InputExc
				[8+ 23 + 2] GRS
				[8+ 23 + 1] Sp
				[8+ 23:23] NormE
				[23-1:0] NormM
			*/
			pipe_2 = {pipe_1[4:0], GRS, Sp, NormE[8:0], NormM[23-1:0]} ;
			/* PIPE 3
				[2*8+2*23+10:2*8+2*23+6] InputExc
				[2*8+2*23+5] GRS
				[2*8+2*23+4] Sp	
				[2*8+2*23+3:8+2*23+3] RoundE
				[8+2*23+2:2*23+2] RoundEP
				[2*23+1:23+1] RoundM
				[23:0] RoundMP
			*/
			pipe_3 = {pipe_2[8+23+7:8+23+1], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]} ;
			/* PIPE 4
				[32+4:5] Z
				[4:0] Flags
			*/				
			pipe_4 = {Z_int[32-1:0], Flags_int[4:0]} ;
		end
	end
		
endmodule



module FPMult_PrepModule (
		clk,
		rst,
		a,
		b,
		Sa,
		Sb,
		Ea,
		Eb,
		Mp,
		InputExc
	);
	
	// Input ports
	input clk ;
	input rst ;
	input [16-1:0] a ;								// Input A, a 32-bit floating point number
	input [16-1:0] b ;								// Input B, a 32-bit floating point number
	
	// Output ports
	output Sa ;										// A's sign
	output Sb ;										// B's sign
	output [8-1:0] Ea ;								// A's exponent
	output [8-1:0] Eb ;								// B's exponent
	output [2*7+1:0] Mp ;							// 7 product
	output [4:0] InputExc ;						// Input numbers are exceptions
	
	// Internal signals							// If signal is high...
	wire ANaN ;										// A is a signalling NaN
	wire BNaN ;										// B is a signalling NaN
	wire AInf ;										// A is infinity
	wire BInf ;										// B is infinity
    wire [7-1:0] Ma;
    wire [7-1:0] Mb;
	
	assign ANaN = &(a[16-2:7]) &  |(a[16-2:7]) ;			// All one 8and not all zero 7 - NaN
	assign BNaN = &(b[16-2:7]) &  |(b[7-1:0]);			// All one 8and not all zero 7 - NaN
	assign AInf = &(a[16-2:7]) & ~|(a[16-2:7]) ;		// All one 8and all zero 7 - Infinity
	assign BInf = &(b[16-2:7]) & ~|(b[16-2:7]) ;		// All one 8and all zero 7 - Infinity
	
	// Check for any exceptions and put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	//assign InputExc = {(ANaN | ANaN | BNaN |BNaN), ANaN, ANaN, BNaN,BNaN} ;
	
	// Take input numbers apart
	assign Sa = a[16-1] ;							// A's sign
	assign Sb = b[16-1] ;							// B's sign
	assign Ea = a[16-2:7];						// Store A's 8in Ea, unless A is an exception
	assign Eb = b[16-2:7];						// Store B's 8in Eb, unless B is an exception	
//    assign Ma = a[7_MSB:7_LSB];
  //  assign Mb = b[7_MSB:7_LSB];
	

	// Actual 7 multiplication occurs here
	//assign Mp = ({4'b0001, a[7-1:0]}*{4'b0001, b[7-1:9]}) ;
	assign Mp = ({1'b1,a[7-1:0]}*{1'b1, b[7-1:0]}) ;

	
    //We multiply part of the 7 here
    //Full 7 of A
    //Bits 7_MUL_SPLIT_MSB:7_MUL_SPLIT_LSB of B
   // wire [`ACTUAL_7-1:0] inp_A;
   // wire [`ACTUAL_7-1:0] inp_B;
   // assign inp_A = {1'b1, Ma};
   // assign inp_B = {{(7-(7_MUL_SPLIT_MSB-7_MUL_SPLIT_LSB+1)){1'b0}}, 1'b1, Mb[7_MUL_SPLIT_MSB:7_MUL_SPLIT_LSB]};
   // DW02_mult #(`ACTUAL_7,`ACTUAL_7) u_mult(.A(inp_A), .B(inp_B), .TC(1'b0), .PRODUCT(Mp));
endmodule


module FPMult_ExecuteModule(
		a,
		b,
		MpC,
		Ea,
		Eb,
		Sa,
		Sb,
		Sp,
		NormE,
		NormM,
		GRS
    );

	// Input ports
	input [7-1:0] a ;
	input [2*8:0] b ;
	input [2*7+1:0] MpC ;
	input [8-1:0] Ea ;						// A's exponent
	input [8-1:0] Eb ;						// B's exponent
	input Sa ;								// A's sign
	input Sb ;								// B's sign
	
	// Output ports
	output Sp ;								// Product sign
	output [8:0] NormE ;													// Normalized exponent
	output [23-1:0] NormM ;												// Normalized 7
	output GRS ;
	
	wire [2*7+1:0] Mp ;
	
	assign Sp = (Sa ^ Sb) ;												// Equal signs give a positive product
	
   // wire [`ACTUAL_7-1:0] inp_a;
   // wire [`ACTUAL_7-1:0] inp_b;
   // assign inp_a = {1'b1, a};
   // assign inp_b = {{(7-7_MUL_SPLIT_LSB){1'b0}}, 1'b0, b};
   // DW02_mult #(`ACTUAL_7,`ACTUAL_7) u_mult(.A(inp_a), .B(inp_b), .TC(1'b0), .PRODUCT(Mp_temp));
   // DW01_add #(2*`ACTUAL_7) u_add(.A(Mp_temp), .B(MpC<<7_MUL_SPLIT_LSB), .CI(1'b0), .SUM(Mp), .CO());

	//assign Mp = (MpC<<(2*8+1)) + ({4'b0001, a[7-1:0]}*{1'b0, b[2*8:0]}) ;
	assign Mp = MpC;


	assign NormM = (Mp[2*7+1] ? Mp[2*7:0] : Mp[2*7-1:0]); 	// Check for overflow
	assign NormE = (Ea + Eb + Mp[2*7+1]);								// If so, increment exponent
	
	assign GRS = ((Mp[7]&(Mp[7+1]))|(|Mp[7-1:0])) ;
	
endmodule

module FPMult_NormalizeModule(
		NormM,
		NormE,
		RoundE,
		RoundEP,
		RoundM,
		RoundMP
    );

	// Input Ports
	input [23-1:0] NormM ;									// Normalized 7
	input [8:0] NormE ;									// Normalized exponent

	// Output Ports
	output [8:0] RoundE ;
	output [8:0] RoundEP ;
	output [23:0] RoundM ;
	output [23:0] RoundMP ; 
	
// 8= 5 
// 8-1 = 4
// NEED to subtract 2^4 -1 = 15

//wire [8-1 : 0] bias;

//assign bias =  ((1<< (8-1)) -1);

	assign RoundE = NormE - 9'd127 ;
	assign RoundEP = NormE - 9'd127 -1 ;
	assign RoundM = NormM ;
	assign RoundMP = NormM ;

endmodule

module FPMult_RoundModule(
		RoundM,
		RoundMP,
		RoundE,
		RoundEP,
		Sp,
		GRS,
		InputExc,
		Z,
		Flags
    );

	// Input Ports
	input [23:0] RoundM ;									// Normalized 7
	input [23:0] RoundMP ;									// Normalized exponent
	input [8:0] RoundE ;									// Normalized 7 + 1
	input [8:0] RoundEP ;									// Normalized 8+ 1
	input Sp ;												// Product sign
	input GRS ;
	input [4:0] InputExc ;
	
	// Output Ports
	output [32-1:0] Z ;										// Final product
	output [4:0] Flags ;
	
	// Internal Signals
	wire [8:0] FinalE ;									// Rounded exponent
	wire [23:0] FinalM;
	wire [23:0] PreShiftM;
	
	assign PreShiftM = GRS ? RoundMP : RoundM ;	// Round up if R and (G or S)
	
	// Post rounding normalization (potential one bit shift> use shifted 7 if there is overflow)
	assign FinalM = (PreShiftM[23] ? {1'b0, PreShiftM[23:1]} : PreShiftM[23:0]) ;
	
	assign FinalE = (PreShiftM[23] ? RoundEP : RoundE) ; // Increment 8if a shift was done
	
	assign Z = {Sp, FinalE[8-1:0], FinalM[14-1:0], 9'b0} ;   // Putting the pieces together
	assign Flags = InputExc[4:0];

endmodule



`timescale 1ns / 1ps
//`define complex_dsp
`define DWIDTH 16
`define AWIDTH 10
`define MEM_SIZE 1024

`define MAT_MUL_SIZE 4
`define MASK_WIDTH 4
`define LOG2_MAT_MUL_SIZE 2

`define NUM_CYCLES_IN_MAC 3
`define MEM_ACCESS_LATENCY 1
`define REG_DATAWIDTH 32
`define REG_ADDRWIDTH 8
`define ADDR_STRIDE_WIDTH 10
`define MAX_BITS_POOL 3
`define EXPONENT 5
`define MANTISSA 10
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/10/2020 11:43:24 PM
// Design Name: 
// Module Name: matmul_4x4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module matmul_4x4_fp_systolic(
 clk,
 reset,
 pe_reset,
 start_mat_mul,
 done_mat_mul,
 address_mat_a,
 address_mat_b,
 address_mat_c,
 address_stride_a,
 address_stride_b,
 address_stride_c,
 a_data,
 b_data,
 a_data_in, //Data values coming in from previous matmul - systolic connections
 b_data_in,
 c_data_in, //Data values coming in from previous matmul - systolic shifting
 c_data_out, //Data values going out to next matmul - systolic shifting
 a_data_out,
 b_data_out,
 a_addr,
 b_addr,
 c_addr,
 c_data_available,
 validity_mask_a_rows,
 validity_mask_a_cols_b_rows,
 validity_mask_b_cols,
 final_mat_mul_size,
 a_loc,
 b_loc
);

 input clk;
 input reset;
 input pe_reset;
 input start_mat_mul;
 output done_mat_mul;
 input [`AWIDTH-1:0] address_mat_a;
 input [`AWIDTH-1:0] address_mat_b;
 input [`AWIDTH-1:0] address_mat_c;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_a;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_b;
 input [`ADDR_STRIDE_WIDTH-1:0] address_stride_c;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_in;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_in;
 input [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_in;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_out;
 output [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_out;
 output [`AWIDTH-1:0] a_addr;
 output [`AWIDTH-1:0] b_addr;
 output [`AWIDTH-1:0] c_addr;
 output c_data_available;
 input [`MASK_WIDTH-1:0] validity_mask_a_rows;
 input [`MASK_WIDTH-1:0] validity_mask_a_cols_b_rows;
 input [`MASK_WIDTH-1:0] validity_mask_b_cols;
//7:0 is okay here. We aren't going to make a matmul larger than 128x128
//In fact, these will get optimized out by the synthesis tool, because
//we hardcode them at the instantiation level.
 input [7:0] final_mat_mul_size;
 input [7:0] a_loc;
 input [7:0] b_loc;

//////////////////////////////////////////////////////////////////////////
// Logic for clock counting and when to assert done
//////////////////////////////////////////////////////////////////////////

reg done_mat_mul;
//This is 7 bits because the expectation is that clock count will be pretty
//small. For large matmuls, this will need to increased to have more bits.
//In general, a systolic multiplier takes 4*N-2+P cycles, where N is the size 
//of the matmul and P is the number of pipleine stages in the MAC block.
reg [7:0] clk_cnt;

//Finding out number of cycles to assert matmul done.
//When we have to save the outputs to accumulators, then we don't need to
//shift out data. So, we can assert done_mat_mul early.
//In the normal case, we have to include the time to shift out the results. 
//Note: the count expression used to contain "4*final_mat_mul_size", but 
//to avoid multiplication, we now use "final_mat_mul_size<<2"
wire [7:0] clk_cnt_for_done;
assign clk_cnt_for_done = 
                          ((final_mat_mul_size<<2) - 2 + `NUM_CYCLES_IN_MAC) ;  

always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    clk_cnt <= 0;
    done_mat_mul <= 0;
  end
  else if (clk_cnt == clk_cnt_for_done) begin
    done_mat_mul <= 1;
    clk_cnt <= clk_cnt + 1;
  end
  else if (done_mat_mul == 0) begin
    clk_cnt <= clk_cnt + 1;
  end    
  else begin
    done_mat_mul <= 0;
    clk_cnt <= clk_cnt + 1;
  end
end


wire [`DWIDTH-1:0] a0_data;
wire [`DWIDTH-1:0] a1_data;
wire [`DWIDTH-1:0] a2_data;
wire [`DWIDTH-1:0] a3_data;
wire [`DWIDTH-1:0] b0_data;
wire [`DWIDTH-1:0] b1_data;
wire [`DWIDTH-1:0] b2_data;
wire [`DWIDTH-1:0] b3_data;
wire [`DWIDTH-1:0] a1_data_delayed_1;
wire [`DWIDTH-1:0] a2_data_delayed_1;
wire [`DWIDTH-1:0] a2_data_delayed_2;
wire [`DWIDTH-1:0] a3_data_delayed_1;
wire [`DWIDTH-1:0] a3_data_delayed_2;
wire [`DWIDTH-1:0] a3_data_delayed_3;
wire [`DWIDTH-1:0] b1_data_delayed_1;
wire [`DWIDTH-1:0] b2_data_delayed_1;
wire [`DWIDTH-1:0] b2_data_delayed_2;
wire [`DWIDTH-1:0] b3_data_delayed_1;
wire [`DWIDTH-1:0] b3_data_delayed_2;
wire [`DWIDTH-1:0] b3_data_delayed_3;

//////////////////////////////////////////////////////////////////////////
// Instantiation of systolic data setup
//////////////////////////////////////////////////////////////////////////
systolic_data_setup_systolic_4x4_fp u_systolic_data_setup_systolic_4x4_fp(
.clk(clk),
.reset(reset),
.start_mat_mul(start_mat_mul),
.a_addr(a_addr),
.b_addr(b_addr),
.address_mat_a(address_mat_a),
.address_mat_b(address_mat_b),
.address_stride_a(address_stride_a),
.address_stride_b(address_stride_b),
.a_data(a_data),
.b_data(b_data),
.clk_cnt(clk_cnt),
.a0_data(a0_data),
.a1_data_delayed_1(a1_data_delayed_1),
.a2_data_delayed_2(a2_data_delayed_2),
.a3_data_delayed_3(a3_data_delayed_3),
.b0_data(b0_data),
.b1_data_delayed_1(b1_data_delayed_1),
.b2_data_delayed_2(b2_data_delayed_2),
.b3_data_delayed_3(b3_data_delayed_3),
.validity_mask_a_rows(validity_mask_a_rows),
.validity_mask_a_cols_b_rows(validity_mask_a_cols_b_rows),
.validity_mask_b_cols(validity_mask_b_cols),
.final_mat_mul_size(final_mat_mul_size),
.a_loc(a_loc),
.b_loc(b_loc)
);


//////////////////////////////////////////////////////////////////////////
// Logic to mux data_in coming from neighboring matmuls
//////////////////////////////////////////////////////////////////////////
wire [`DWIDTH-1:0] a0;
wire [`DWIDTH-1:0] a1;
wire [`DWIDTH-1:0] a2;
wire [`DWIDTH-1:0] a3;
wire [`DWIDTH-1:0] b0;
wire [`DWIDTH-1:0] b1;
wire [`DWIDTH-1:0] b2;
wire [`DWIDTH-1:0] b3;

wire [`DWIDTH-1:0] a0_data_in;
wire [`DWIDTH-1:0] a1_data_in;
wire [`DWIDTH-1:0] a2_data_in;
wire [`DWIDTH-1:0] a3_data_in;
assign a0_data_in = a_data_in[`DWIDTH-1:0];
assign a1_data_in = a_data_in[2*`DWIDTH-1:`DWIDTH];
assign a2_data_in = a_data_in[3*`DWIDTH-1:2*`DWIDTH];
assign a3_data_in = a_data_in[4*`DWIDTH-1:3*`DWIDTH];

wire [`DWIDTH-1:0] b0_data_in;
wire [`DWIDTH-1:0] b1_data_in;
wire [`DWIDTH-1:0] b2_data_in;
wire [`DWIDTH-1:0] b3_data_in;
assign b0_data_in = b_data_in[`DWIDTH-1:0];
assign b1_data_in = b_data_in[2*`DWIDTH-1:`DWIDTH];
assign b2_data_in = b_data_in[3*`DWIDTH-1:2*`DWIDTH];
assign b3_data_in = b_data_in[4*`DWIDTH-1:3*`DWIDTH];

//If b_loc is 0, that means this matmul block is on the top-row of the
//final large matmul. In that case, b will take inputs from mem.
//If b_loc != 0, that means this matmul block is not on the top-row of the
//final large matmul. In that case, b will take inputs from the matmul on top
//of this one.
assign a0 = (b_loc==0) ? a0_data           : a0_data_in;
assign a1 = (b_loc==0) ? a1_data_delayed_1 : a1_data_in;
assign a2 = (b_loc==0) ? a2_data_delayed_2 : a2_data_in;
assign a3 = (b_loc==0) ? a3_data_delayed_3 : a3_data_in;

//If a_loc is 0, that means this matmul block is on the left-col of the
//final large matmul. In that case, a will take inputs from mem.
//If a_loc != 0, that means this matmul block is not on the left-col of the
//final large matmul. In that case, a will take inputs from the matmul on left
//of this one.
assign b0 = (a_loc==0) ? b0_data           : b0_data_in;
assign b1 = (a_loc==0) ? b1_data_delayed_1 : b1_data_in;
assign b2 = (a_loc==0) ? b2_data_delayed_2 : b2_data_in;
assign b3 = (a_loc==0) ? b3_data_delayed_3 : b3_data_in;


wire [`DWIDTH-1:0] matrixC00;
wire [`DWIDTH-1:0] matrixC01;
wire [`DWIDTH-1:0] matrixC02;
wire [`DWIDTH-1:0] matrixC03;
wire [`DWIDTH-1:0] matrixC10;
wire [`DWIDTH-1:0] matrixC11;
wire [`DWIDTH-1:0] matrixC12;
wire [`DWIDTH-1:0] matrixC13;
wire [`DWIDTH-1:0] matrixC20;
wire [`DWIDTH-1:0] matrixC21;
wire [`DWIDTH-1:0] matrixC22;
wire [`DWIDTH-1:0] matrixC23;
wire [`DWIDTH-1:0] matrixC30;
wire [`DWIDTH-1:0] matrixC31;
wire [`DWIDTH-1:0] matrixC32;
wire [`DWIDTH-1:0] matrixC33;


//////////////////////////////////////////////////////////////////////////
// Instantiation of the output logic
//////////////////////////////////////////////////////////////////////////
output_logic_systolic_4x4_fp u_output_logic_systolic_4x4_fp(
.clk(clk),
.reset(reset),
.start_mat_mul(start_mat_mul),
.done_mat_mul(done_mat_mul),
.address_mat_c(address_mat_c),
.address_stride_c(address_stride_c),
.c_data_out(c_data_out),
.c_data_in(c_data_in),
.c_addr(c_addr),
.c_data_available(c_data_available),
.clk_cnt(clk_cnt),
.final_mat_mul_size(final_mat_mul_size),
.matrixC00(matrixC00),
.matrixC01(matrixC01),
.matrixC02(matrixC02),
.matrixC03(matrixC03),
.matrixC10(matrixC10),
.matrixC11(matrixC11),
.matrixC12(matrixC12),
.matrixC13(matrixC13),
.matrixC20(matrixC20),
.matrixC21(matrixC21),
.matrixC22(matrixC22),
.matrixC23(matrixC23),
.matrixC30(matrixC30),
.matrixC31(matrixC31),
.matrixC32(matrixC32),
.matrixC33(matrixC33)
);

//////////////////////////////////////////////////////////////////////////
// Instantiations of the actual PEs
//////////////////////////////////////////////////////////////////////////
systolic_pe_matrix_systolic_4x4_fp u_systolic_pe_matrix_systolic_4x4_fp(
.reset(reset),
.clk(clk),
.pe_reset(pe_reset),
.start_mat_mul(start_mat_mul),
.a0(a0), 
.a1(a1), 
.a2(a2), 
.a3(a3),
.b0(b0), 
.b1(b1), 
.b2(b2), 
.b3(b3),
.matrixC00(matrixC00),
.matrixC01(matrixC01),
.matrixC02(matrixC02),
.matrixC03(matrixC03),
.matrixC10(matrixC10),
.matrixC11(matrixC11),
.matrixC12(matrixC12),
.matrixC13(matrixC13),
.matrixC20(matrixC20),
.matrixC21(matrixC21),
.matrixC22(matrixC22),
.matrixC23(matrixC23),
.matrixC30(matrixC30),
.matrixC31(matrixC31),
.matrixC32(matrixC32),
.matrixC33(matrixC33),
.a_data_out(a_data_out),
.b_data_out(b_data_out)
);

endmodule

//////////////////////////////////////////////////////////////////////////
// Output logic
//////////////////////////////////////////////////////////////////////////
module output_logic_systolic_4x4_fp(
clk,
reset,
start_mat_mul,
done_mat_mul,
address_mat_c,
address_stride_c,
c_data_in,
c_data_out, //Data values going out to next matmul - systolic shifting
c_addr,
c_data_available,
clk_cnt,
final_mat_mul_size,
matrixC00,
matrixC01,
matrixC02,
matrixC03,
matrixC10,
matrixC11,
matrixC12,
matrixC13,
matrixC20,
matrixC21,
matrixC22,
matrixC23,
matrixC30,
matrixC31,
matrixC32,
matrixC33
);

input clk;
input reset;
input start_mat_mul;
input done_mat_mul;
input [`AWIDTH-1:0] address_mat_c;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_c;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_in;
output [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out;
output [`AWIDTH-1:0] c_addr;
output c_data_available;
input [7:0] clk_cnt;
//output row_latch_en;
input [7:0] final_mat_mul_size;
input [`DWIDTH-1:0] matrixC00;
input [`DWIDTH-1:0] matrixC01;
input [`DWIDTH-1:0] matrixC02;
input [`DWIDTH-1:0] matrixC03;
input [`DWIDTH-1:0] matrixC10;
input [`DWIDTH-1:0] matrixC11;
input [`DWIDTH-1:0] matrixC12;
input [`DWIDTH-1:0] matrixC13;
input [`DWIDTH-1:0] matrixC20;
input [`DWIDTH-1:0] matrixC21;
input [`DWIDTH-1:0] matrixC22;
input [`DWIDTH-1:0] matrixC23;
input [`DWIDTH-1:0] matrixC30;
input [`DWIDTH-1:0] matrixC31;
input [`DWIDTH-1:0] matrixC32;
input [`DWIDTH-1:0] matrixC33;

wire row_latch_en;

//////////////////////////////////////////////////////////////////////////
// Logic to capture matrix C data from the PEs and shift it out
//////////////////////////////////////////////////////////////////////////

//assign row_latch_en = (clk_cnt==(`MAT_MUL_SIZE + (a_loc+b_loc) * `BB_MAT_MUL_SIZE + 10 +  `NUM_CYCLES_IN_MAC - 1));
//Writing the line above to avoid multiplication:
//assign row_latch_en = (clk_cnt==(`MAT_MUL_SIZE + ((a_loc+b_loc) << `LOG2_MAT_MUL_SIZE) + 10 +  `NUM_CYCLES_IN_MAC - 1));
//Fixing bug. The line above is inaccurate. Using the line below. 
//TODO: This line needs to be fixed to include a_loc and b_loc ie. when final_mat_mul_size is different from `MAT_MUL_SIZE
assign row_latch_en =  
                       //((clk_cnt == ((`MAT_MUL_SIZE<<2) - `MAT_MUL_SIZE -2 +`NUM_CYCLES_IN_MAC)));
                       ((clk_cnt == ((final_mat_mul_size<<2) - final_mat_mul_size -1 +`NUM_CYCLES_IN_MAC)));

reg c_data_available;
reg [`AWIDTH-1:0] c_addr;
reg start_capturing_c_data;
integer counter;
reg [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out;
reg [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out_1;
reg [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out_2;
reg [`MAT_MUL_SIZE*`DWIDTH-1:0] c_data_out_3;

wire [`MAT_MUL_SIZE*`DWIDTH-1:0] col0;
wire [`MAT_MUL_SIZE*`DWIDTH-1:0] col1;
wire [`MAT_MUL_SIZE*`DWIDTH-1:0] col2;
wire [`MAT_MUL_SIZE*`DWIDTH-1:0] col3;
assign col0 = {matrixC30, matrixC20, matrixC10, matrixC00};
assign col1 = {matrixC31, matrixC21, matrixC11, matrixC01};
assign col2 = {matrixC32, matrixC22, matrixC12, matrixC02};
assign col3 = {matrixC33, matrixC23, matrixC13, matrixC03};

//If save_output_to_accum is asserted, that means we are not intending to shift
//out the outputs, because the outputs are still partial sums. 
wire condition_to_start_shifting_output;
assign condition_to_start_shifting_output = 
                          row_latch_en ;  

//For larger matmuls, this logic will have more entries in the case statement
always @(posedge clk) begin
  if (reset | ~start_mat_mul) begin
    start_capturing_c_data <= 1'b0;
    c_data_available <= 1'b0;
    c_addr <= address_mat_c+address_stride_c;
    c_data_out <= 0;
    counter <= 0;
    c_data_out_1 <= 0; 
    c_data_out_2 <= 0; 
    c_data_out_3 <= 0; 
  end
  else if (condition_to_start_shifting_output) begin
    start_capturing_c_data <= 1'b1;
    c_data_available <= 1'b1;
    c_addr <= c_addr - address_stride_c;
    c_data_out <= col0; 
    c_data_out_1 <= col1; 
    c_data_out_2 <= col2; 
    c_data_out_3 <= col3; 
    counter <= counter + 1;
  end 
  else if (done_mat_mul) begin
    start_capturing_c_data <= 1'b0;
    c_data_available <= 1'b0;
    c_addr <= address_mat_c+address_stride_c;
    c_data_out <= 0;
    c_data_out_1 <= 0;
    c_data_out_2 <= 0;
    c_data_out_3 <= 0;
  end 
  else if (counter >= `MAT_MUL_SIZE) begin
    c_addr <= c_addr - address_stride_c;
    c_data_out <= c_data_out_1;
    c_data_out_1 <= c_data_out_2;
    c_data_out_2 <= c_data_out_3;
    c_data_out_3 <= c_data_in;
  end
  else if (start_capturing_c_data) begin
    c_data_available <= 1'b1;
    c_addr <= c_addr - address_stride_c;
    counter <= counter + 1;
    c_data_out <= c_data_out_1;
    c_data_out_1 <= c_data_out_2;
    c_data_out_2 <= c_data_out_3;
    c_data_out_3 <= c_data_in;
  end
end

endmodule

//////////////////////////////////////////////////////////////////////////
// Systolic data setup
//////////////////////////////////////////////////////////////////////////
module systolic_data_setup_systolic_4x4_fp(
clk,
reset,
start_mat_mul,
a_addr,
b_addr,
address_mat_a,
address_mat_b,
address_stride_a,
address_stride_b,
a_data,
b_data,
clk_cnt,
a0_data,
a1_data_delayed_1,
a2_data_delayed_2,
a3_data_delayed_3,
b0_data,
b1_data_delayed_1,
b2_data_delayed_2,
b3_data_delayed_3,
validity_mask_a_rows,
validity_mask_a_cols_b_rows,
validity_mask_b_cols,
final_mat_mul_size,
a_loc,
b_loc
);

input clk;
input reset;
input start_mat_mul;
output [`AWIDTH-1:0] a_addr;
output [`AWIDTH-1:0] b_addr;
input [`AWIDTH-1:0] address_mat_a;
input [`AWIDTH-1:0] address_mat_b;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_a;
input [`ADDR_STRIDE_WIDTH-1:0] address_stride_b;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data;
input [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data;
input [7:0] clk_cnt;
output [`DWIDTH-1:0] a0_data;
output [`DWIDTH-1:0] a1_data_delayed_1;
output [`DWIDTH-1:0] a2_data_delayed_2;
output [`DWIDTH-1:0] a3_data_delayed_3;
output [`DWIDTH-1:0] b0_data;
output [`DWIDTH-1:0] b1_data_delayed_1;
output [`DWIDTH-1:0] b2_data_delayed_2;
output [`DWIDTH-1:0] b3_data_delayed_3;
input [`MASK_WIDTH-1:0] validity_mask_a_rows;
input [`MASK_WIDTH-1:0] validity_mask_a_cols_b_rows;
input [`MASK_WIDTH-1:0] validity_mask_b_cols;
input [7:0] final_mat_mul_size;
input [7:0] a_loc;
input [7:0] b_loc;

wire [`DWIDTH-1:0] a0_data;
wire [`DWIDTH-1:0] a1_data;
wire [`DWIDTH-1:0] a2_data;
wire [`DWIDTH-1:0] a3_data;
wire [`DWIDTH-1:0] b0_data;
wire [`DWIDTH-1:0] b1_data;
wire [`DWIDTH-1:0] b2_data;
wire [`DWIDTH-1:0] b3_data;

//////////////////////////////////////////////////////////////////////////
// Logic to generate addresses to BRAM A
//////////////////////////////////////////////////////////////////////////
reg [`AWIDTH-1:0] a_addr;
reg a_mem_access; //flag that tells whether the matmul is trying to access memory or not

always @(posedge clk) begin
  //else if (clk_cnt >= a_loc*`MAT_MUL_SIZE+final_mat_mul_size) begin
  //Writing the line above to avoid multiplication:
  if ((reset || ~start_mat_mul) || (clk_cnt >= (a_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
      a_addr <= address_mat_a-address_stride_a;
    a_mem_access <= 0;
  end

  //else if ((clk_cnt >= a_loc*`MAT_MUL_SIZE) && (clk_cnt < a_loc*`MAT_MUL_SIZE+final_mat_mul_size)) begin
  //Writing the line above to avoid multiplication:
  else if ((clk_cnt >= (a_loc<<`LOG2_MAT_MUL_SIZE)) && (clk_cnt < (a_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
      a_addr <= a_addr + address_stride_a;
    a_mem_access <= 1;
  end
end  

//////////////////////////////////////////////////////////////////////////
// Logic to generate valid signals for data coming from BRAM A
//////////////////////////////////////////////////////////////////////////
reg [7:0] a_mem_access_counter;
always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    a_mem_access_counter <= 0;
  end
  else if (a_mem_access == 1) begin
    a_mem_access_counter <= a_mem_access_counter + 1;  

  end
  else begin
    a_mem_access_counter <= 0;
  end
end

wire a_data_valid; //flag that tells whether the data from memory is valid
assign a_data_valid = 
       ((validity_mask_a_cols_b_rows[0]==1'b0 && a_mem_access_counter==1) ||
        (validity_mask_a_cols_b_rows[1]==1'b0 && a_mem_access_counter==2) ||
        (validity_mask_a_cols_b_rows[2]==1'b0 && a_mem_access_counter==3) ||
        (validity_mask_a_cols_b_rows[3]==1'b0 && a_mem_access_counter==4)) ?
        1'b0 : (a_mem_access_counter >= `MEM_ACCESS_LATENCY);

//////////////////////////////////////////////////////////////////////////
// Logic to delay certain parts of the data received from BRAM A (systolic data setup)
//////////////////////////////////////////////////////////////////////////
//Slice data into chunks and qualify it with whether it is valid or not
assign a0_data = a_data[`DWIDTH-1:0] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[0]}};
assign a1_data = a_data[2*`DWIDTH-1:`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[1]}};
assign a2_data = a_data[3*`DWIDTH-1:2*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[2]}};
assign a3_data = a_data[4*`DWIDTH-1:3*`DWIDTH] & {`DWIDTH{a_data_valid}} & {`DWIDTH{validity_mask_a_rows[3]}};

//For larger matmuls, more such delaying flops will be needed
reg [`DWIDTH-1:0] a1_data_delayed_1;
reg [`DWIDTH-1:0] a2_data_delayed_1;
reg [`DWIDTH-1:0] a2_data_delayed_2;
reg [`DWIDTH-1:0] a3_data_delayed_1;
reg [`DWIDTH-1:0] a3_data_delayed_2;
reg [`DWIDTH-1:0] a3_data_delayed_3;
always @(posedge clk) begin
  if (reset || ~start_mat_mul || clk_cnt==0) begin
    a1_data_delayed_1 <= 0;
    a2_data_delayed_1 <= 0;
    a2_data_delayed_2 <= 0;
    a3_data_delayed_1 <= 0;
    a3_data_delayed_2 <= 0;
    a3_data_delayed_3 <= 0;
  end
  else begin
    a1_data_delayed_1 <= a1_data;
    a2_data_delayed_1 <= a2_data;
    a2_data_delayed_2 <= a2_data_delayed_1;
    a3_data_delayed_1 <= a3_data;
    a3_data_delayed_2 <= a3_data_delayed_1;
    a3_data_delayed_3 <= a3_data_delayed_2;
  end
end

//////////////////////////////////////////////////////////////////////////
// Logic to generate addresses to BRAM B
//////////////////////////////////////////////////////////////////////////
reg [`AWIDTH-1:0] b_addr;
reg b_mem_access; //flag that tells whether the matmul is trying to access memory or not

always @(posedge clk) begin
  //else if (clk_cnt >= b_loc*`MAT_MUL_SIZE+final_mat_mul_size) begin
  //Writing the line above to avoid multiplication:
  if ((reset || ~start_mat_mul) || (clk_cnt >= (b_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
      b_addr <= address_mat_b - address_stride_b;
    b_mem_access <= 0;
  end
  //else if ((clk_cnt >= b_loc*`MAT_MUL_SIZE) && (clk_cnt < b_loc*`MAT_MUL_SIZE+final_mat_mul_size)) begin
  //Writing the line above to avoid multiplication:
  else if ((clk_cnt >= (b_loc<<`LOG2_MAT_MUL_SIZE)) && (clk_cnt < (b_loc<<`LOG2_MAT_MUL_SIZE)+final_mat_mul_size)) begin
      b_addr <= b_addr + address_stride_b;
    b_mem_access <= 1;
  end
end  

//////////////////////////////////////////////////////////////////////////
// Logic to generate valid signals for data coming from BRAM B
//////////////////////////////////////////////////////////////////////////
reg [7:0] b_mem_access_counter;
always @(posedge clk) begin
  if (reset || ~start_mat_mul) begin
    b_mem_access_counter <= 0;
  end
  else if (b_mem_access == 1) begin
    b_mem_access_counter <= b_mem_access_counter + 1;  
  end
  else begin
    b_mem_access_counter <= 0;
  end
end

wire b_data_valid; //flag that tells whether the data from memory is valid
assign b_data_valid = 
       ((validity_mask_a_cols_b_rows[0]==1'b0 && b_mem_access_counter==1) ||
        (validity_mask_a_cols_b_rows[1]==1'b0 && b_mem_access_counter==2) ||
        (validity_mask_a_cols_b_rows[2]==1'b0 && b_mem_access_counter==3) ||
        (validity_mask_a_cols_b_rows[3]==1'b0 && b_mem_access_counter==4)) ?
        1'b0 : (b_mem_access_counter >= `MEM_ACCESS_LATENCY);


//////////////////////////////////////////////////////////////////////////
// Logic to delay certain parts of the data received from BRAM B (systolic data setup)
//////////////////////////////////////////////////////////////////////////
//Slice data into chunks and qualify it with whether it is valid or not
assign b0_data = b_data[`DWIDTH-1:0] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[0]}};
assign b1_data = b_data[2*`DWIDTH-1:`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[1]}};
assign b2_data = b_data[3*`DWIDTH-1:2*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[2]}};
assign b3_data = b_data[4*`DWIDTH-1:3*`DWIDTH] & {`DWIDTH{b_data_valid}} & {`DWIDTH{validity_mask_b_cols[3]}};

//For larger matmuls, more such delaying flops will be needed
reg [`DWIDTH-1:0] b1_data_delayed_1;
reg [`DWIDTH-1:0] b2_data_delayed_1;
reg [`DWIDTH-1:0] b2_data_delayed_2;
reg [`DWIDTH-1:0] b3_data_delayed_1;
reg [`DWIDTH-1:0] b3_data_delayed_2;
reg [`DWIDTH-1:0] b3_data_delayed_3;
always @(posedge clk) begin
  if (reset || ~start_mat_mul || clk_cnt==0) begin
    b1_data_delayed_1 <= 0;
    b2_data_delayed_1 <= 0;
    b2_data_delayed_2 <= 0;
    b3_data_delayed_1 <= 0;
    b3_data_delayed_2 <= 0;
    b3_data_delayed_3 <= 0;
  end
  else begin
    b1_data_delayed_1 <= b1_data;
    b2_data_delayed_1 <= b2_data;
    b2_data_delayed_2 <= b2_data_delayed_1;
    b3_data_delayed_1 <= b3_data;
    b3_data_delayed_2 <= b3_data_delayed_1;
    b3_data_delayed_3 <= b3_data_delayed_2;
  end
end


endmodule



//////////////////////////////////////////////////////////////////////////
// Systolically connected PEs
//////////////////////////////////////////////////////////////////////////
module systolic_pe_matrix_systolic_4x4_fp(
reset,
clk,
pe_reset,
start_mat_mul,
a0, a1, a2, a3,
b0, b1, b2, b3,
matrixC00,
matrixC01,
matrixC02,
matrixC03,
matrixC10,
matrixC11,
matrixC12,
matrixC13,
matrixC20,
matrixC21,
matrixC22,
matrixC23,
matrixC30,
matrixC31,
matrixC32,
matrixC33,
a_data_out,
b_data_out
);

input clk;
input reset;
input pe_reset;
input start_mat_mul;
input [`DWIDTH-1:0] a0;
input [`DWIDTH-1:0] a1;
input [`DWIDTH-1:0] a2;
input [`DWIDTH-1:0] a3;
input [`DWIDTH-1:0] b0;
input [`DWIDTH-1:0] b1;
input [`DWIDTH-1:0] b2;
input [`DWIDTH-1:0] b3;
output [`DWIDTH-1:0] matrixC00;
output [`DWIDTH-1:0] matrixC01;
output [`DWIDTH-1:0] matrixC02;
output [`DWIDTH-1:0] matrixC03;
output [`DWIDTH-1:0] matrixC10;
output [`DWIDTH-1:0] matrixC11;
output [`DWIDTH-1:0] matrixC12;
output [`DWIDTH-1:0] matrixC13;
output [`DWIDTH-1:0] matrixC20;
output [`DWIDTH-1:0] matrixC21;
output [`DWIDTH-1:0] matrixC22;
output [`DWIDTH-1:0] matrixC23;
output [`DWIDTH-1:0] matrixC30;
output [`DWIDTH-1:0] matrixC31;
output [`DWIDTH-1:0] matrixC32;
output [`DWIDTH-1:0] matrixC33;
output [`MAT_MUL_SIZE*`DWIDTH-1:0] a_data_out;
output [`MAT_MUL_SIZE*`DWIDTH-1:0] b_data_out;

wire [`DWIDTH-1:0] a00to01, a01to02, a02to03, a03to04;
wire [`DWIDTH-1:0] a10to11, a11to12, a12to13, a13to14;
wire [`DWIDTH-1:0] a20to21, a21to22, a22to23, a23to24;
wire [`DWIDTH-1:0] a30to31, a31to32, a32to33, a33to34;

wire [`DWIDTH-1:0] b00to10, b10to20, b20to30, b30to40; 
wire [`DWIDTH-1:0] b01to11, b11to21, b21to31, b31to41;
wire [`DWIDTH-1:0] b02to12, b12to22, b22to32, b32to42;
wire [`DWIDTH-1:0] b03to13, b13to23, b23to33, b33to43;

wire effective_rst;
assign effective_rst = reset | pe_reset;

 processing_element_systolic_4x4_fp pe00(.reset(effective_rst), .clk(clk),  .in_a(a0),      .in_b(b0),  .out_a(a00to01), .out_b(b00to10), .out_c(matrixC00));
 processing_element_systolic_4x4_fp pe01(.reset(effective_rst), .clk(clk),  .in_a(a00to01), .in_b(b1),  .out_a(a01to02), .out_b(b01to11), .out_c(matrixC01));
 processing_element_systolic_4x4_fp pe02(.reset(effective_rst), .clk(clk),  .in_a(a01to02), .in_b(b2),  .out_a(a02to03), .out_b(b02to12), .out_c(matrixC02));
 processing_element_systolic_4x4_fp pe03(.reset(effective_rst), .clk(clk),  .in_a(a02to03), .in_b(b3),  .out_a(a03to04), .out_b(b03to13), .out_c(matrixC03));

 processing_element_systolic_4x4_fp pe10(.reset(effective_rst), .clk(clk),  .in_a(a1),      .in_b(b00to10), .out_a(a10to11), .out_b(b10to20), .out_c(matrixC10));
 processing_element_systolic_4x4_fp pe11(.reset(effective_rst), .clk(clk),  .in_a(a10to11), .in_b(b01to11), .out_a(a11to12), .out_b(b11to21), .out_c(matrixC11));
 processing_element_systolic_4x4_fp pe12(.reset(effective_rst), .clk(clk),  .in_a(a11to12), .in_b(b02to12), .out_a(a12to13), .out_b(b12to22), .out_c(matrixC12));
 processing_element_systolic_4x4_fp pe13(.reset(effective_rst), .clk(clk),  .in_a(a12to13), .in_b(b03to13), .out_a(a13to14), .out_b(b13to23), .out_c(matrixC13));

 processing_element_systolic_4x4_fp pe20(.reset(effective_rst), .clk(clk),  .in_a(a2),      .in_b(b10to20), .out_a(a20to21), .out_b(b20to30), .out_c(matrixC20));
 processing_element_systolic_4x4_fp pe21(.reset(effective_rst), .clk(clk),  .in_a(a20to21), .in_b(b11to21), .out_a(a21to22), .out_b(b21to31), .out_c(matrixC21));
 processing_element_systolic_4x4_fp pe22(.reset(effective_rst), .clk(clk),  .in_a(a21to22), .in_b(b12to22), .out_a(a22to23), .out_b(b22to32), .out_c(matrixC22));
 processing_element_systolic_4x4_fp pe23(.reset(effective_rst), .clk(clk),  .in_a(a22to23), .in_b(b13to23), .out_a(a23to24), .out_b(b23to33), .out_c(matrixC23));

 processing_element_systolic_4x4_fp pe30(.reset(effective_rst), .clk(clk),  .in_a(a3),      .in_b(b20to30), .out_a(a30to31), .out_b(b30to40), .out_c(matrixC30));
 processing_element_systolic_4x4_fp pe31(.reset(effective_rst), .clk(clk),  .in_a(a30to31), .in_b(b21to31), .out_a(a31to32), .out_b(b31to41), .out_c(matrixC31));
 processing_element_systolic_4x4_fp pe32(.reset(effective_rst), .clk(clk),  .in_a(a31to32), .in_b(b22to32), .out_a(a32to33), .out_b(b32to42), .out_c(matrixC32));
 processing_element_systolic_4x4_fp pe33(.reset(effective_rst), .clk(clk),  .in_a(a32to33), .in_b(b23to33), .out_a(a33to34), .out_b(b33to43), .out_c(matrixC33));

assign a_data_out = {a33to34,a23to24,a13to14,a03to04};
assign b_data_out = {b33to43,b32to42,b31to41,b30to40};

endmodule



//////////////////////////////////////////////////////////////////////////
// Definition of a processing element (basically a MAC)
//////////////////////////////////////////////////////////////////////////
module  processing_element_systolic_4x4_fp(
 reset, 
 clk, 
 in_a,
 in_b, 
 out_a, 
 out_b, 
 out_c
 );

 input reset;
 input clk;
 input  [`DWIDTH-1:0] in_a;
 input  [`DWIDTH-1:0] in_b;
 output [`DWIDTH-1:0] out_a;
 output [`DWIDTH-1:0] out_b;
 output [`DWIDTH-1:0] out_c;  //reduced precision

 reg [`DWIDTH-1:0] out_a;
 reg [`DWIDTH-1:0] out_b;
 wire [`DWIDTH-1:0] out_c;

 wire [`DWIDTH-1:0] out_mac;

 assign out_c = out_mac;

 `ifdef complex_dsp
 mac_fp u_mac(.a(in_a), .b(in_b), .out(out_mac), .reset(reset), .clk(clk));
 `else
 seq_mac_systolic_4x4_fp u_mac(.a(in_a), .b(in_b), .out(out_mac), .reset(reset), .clk(clk));
 `endif

 always @(posedge clk)begin
    if(reset) begin
      out_a<=0;
      out_b<=0;
    end
    else begin  
      out_a<=in_a;
      out_b<=in_b;
    end
 end
 
endmodule

//////////////////////////////////////////////////////////////////////////
// Multiply-and-accumulate (MAC) block
//////////////////////////////////////////////////////////////////////////
//module seq_mac_systolic_4x4_fp(a, b, out, reset, clk);
//input [`DWIDTH-1:0] a;
//input [`DWIDTH-1:0] b;
//input reset;
//input clk;
//output [`DWIDTH-1:0] out;
//
//reg [2*`DWIDTH-1:0] out_temp;
//wire [`DWIDTH-1:0] mul_out;
//wire [2*`DWIDTH-1:0] add_out;
//
//reg [`DWIDTH-1:0] a_flopped;
//reg [`DWIDTH-1:0] b_flopped;
//
//wire [2*`DWIDTH-1:0] mul_out_temp;
//reg [2*`DWIDTH-1:0] mul_out_temp_reg;
//
//always @(posedge clk) begin
//  if (reset) begin
//    a_flopped <= 0;
//    b_flopped <= 0;
//  end else begin
//    a_flopped <= a;
//    b_flopped <= b;
//  end
//end
//
////assign mul_out = a * b;
//qmult_systolic_4x4_fp mult_u1(.i_multiplicand(a_flopped), .i_multiplier(b_flopped), .o_result(mul_out_temp));
//
//always @(posedge clk) begin
//  if (reset) begin
//    mul_out_temp_reg <= 0;
//  end else begin
//    mul_out_temp_reg <= mul_out_temp;
//  end
//end
//
////we just truncate the higher bits of the product
////assign add_out = mul_out + out;
//qadd_systolic_4x4_fp add_u1(.a(out_temp), .b(mul_out_temp_reg), .c(add_out));
//
//always @(posedge clk) begin
//  if (reset) begin
//    out_temp <= 0;
//  end else begin
//    out_temp <= add_out;
//  end
//end
//
////down cast the result
//assign out = 
//    (out_temp[2*`DWIDTH-1] == 0) ?  //positive number
//        (
//           (|(out_temp[2*`DWIDTH-2 : `DWIDTH-1])) ?  //is any bit from 14:7 is 1, that means overlfow
//             {out_temp[2*`DWIDTH-1] , {(`DWIDTH-1){1'b1}}} : //sign bit and then all 1s
//             {out_temp[2*`DWIDTH-1] , out_temp[`DWIDTH-2:0]} 
//        )
//        : //negative number
//        (
//           (|(out_temp[2*`DWIDTH-2 : `DWIDTH-1])) ?  //is any bit from 14:7 is 0, that means overlfow
//             {out_temp[2*`DWIDTH-1] , out_temp[`DWIDTH-2:0]} :
//             {out_temp[2*`DWIDTH-1] , {(`DWIDTH-1){1'b0}}} //sign bit and then all 0s
//        );
//
//endmodule
//
//module qmult_systolic_4x4_fp(i_multiplicand,i_multiplier,o_result);
//input [`DWIDTH-1:0] i_multiplicand;
//input [`DWIDTH-1:0] i_multiplier;
//output [2*`DWIDTH-1:0] o_result;
//
//assign o_result = i_multiplicand * i_multiplier;
////DW02_mult #(`DWIDTH,`DWIDTH) u_mult(.A(i_multiplicand), .B(i_multiplier), .TC(1'b1), .PRODUCT(o_result));
//
//endmodule
//
//module qadd_systolic_4x4_fp(a,b,c);
//input [2*`DWIDTH-1:0] a;
//input [2*`DWIDTH-1:0] b;
//output [2*`DWIDTH-1:0] c;
//
//assign c = a + b;
////DW01_add #(`DWIDTH) u_add(.A(a), .B(b), .CI(1'b0), .SUM(c), .CO());
//endmodule

`ifndef complex_dsp

//////////////////////////////////////////////////////////////////////////
// Multiply-and-accumulate (MAC) block
//////////////////////////////////////////////////////////////////////////
module seq_mac_systolic_4x4_fp(a, b, out, reset, clk);
input [`DWIDTH-1:0] a;
input [`DWIDTH-1:0] b;
input reset;
input clk;
output [`DWIDTH-1:0] out;

reg [2*`DWIDTH-1:0] out_temp;
wire [2*`DWIDTH-1:0] mul_out;
wire [2*`DWIDTH-1:0] add_out;

reg [`DWIDTH-1:0] a_flopped;
reg [`DWIDTH-1:0] b_flopped;

wire [2*`DWIDTH-1:0] mul_out_temp;
reg [2*`DWIDTH-1:0] mul_out_temp_reg;

always @(posedge clk) begin
  if (reset) begin
    a_flopped <= 0;
    b_flopped <= 0;
  end else begin
    a_flopped <= a;
    b_flopped <= b;
  end
end

//assign mul_out = a * b;
qmult_systolic_4x4_fp mult_u1(.clk(clk), .rst(reset), .i_multiplicand(a_flopped), .i_multiplier(b_flopped), .o_result(mul_out_temp));

always @(posedge clk) begin
  if (reset) begin
    mul_out_temp_reg <= 0;
  end else begin
    mul_out_temp_reg <= mul_out_temp;
  end
end

assign mul_out = mul_out_temp_reg;

qadd_systolic_4x4_fp add_u1(.clk(clk), .rst(reset), .a(out_temp), .b(mul_out), .c(add_out));

always @(posedge clk) begin
  if (reset) begin
    out_temp <= 0;
  end else begin
    out_temp <= add_out;
  end
end

//fp32 to fp16 conversion
wire [15:0] fpadd_16_result;
fp32_to_fp16_systolic_4x4_fp u_32to16 (.a(out_temp), .b(out));

endmodule


//////////////////////////////////////////////////////////////////////////
// Multiplier
//////////////////////////////////////////////////////////////////////////
module qmult_systolic_4x4_fp(clk,rst,i_multiplicand,i_multiplier,o_result);
input clk;
input rst;
input [`DWIDTH-1:0] i_multiplicand;
input [`DWIDTH-1:0] i_multiplier;
output [2*`DWIDTH-1:0] o_result;

wire FPMult_16_systolic_4x4_fp_clk_NC;
wire FPMult_16_systolic_4x4_fp_rst_NC;
wire [15:0] FPMult_16_systolic_4x4_fp_result;
wire [4:0] FPMult_16_systolic_4x4_fp_flags;

FPMult_16_systolic_4x4_fp u_FPMult_16_systolic_4x4_fp(
   .clk(clk),
   .rst(rst),
   .a(i_multiplicand[15:0]),
   .b(i_multiplier[15:0]),
   .result(FPMult_16_systolic_4x4_fp_result),
   .flags(FPMult_16_systolic_4x4_fp_flags)
 );

//Convert fp16 to fp32
fp16_to_fp32_systolic_4x4_fp u_16to32 (.a(FPMult_16_systolic_4x4_fp_result), .b(o_result));

endmodule


//////////////////////////////////////////////////////////////////////////
// Adder
//////////////////////////////////////////////////////////////////////////
module qadd_systolic_4x4_fp(clk,rst,a,b,c);
input clk;
input rst;
input [2*`DWIDTH-1:0] a;
input [2*`DWIDTH-1:0] b;
output [2*`DWIDTH-1:0] c;

wire fpadd_32_clk_NC;
wire fpadd_32_rst_NC;
wire [4:0] fpadd_32_flags;

FPAddSub_single_systolic_4x4_fp u_fpaddsub_32(
  .clk(clk),
  .rst(rst),
  .a(a),
  .b(b),
  .operation(1'b0), 
  .result(c),
  .flags(fpadd_32_flags));

endmodule
`endif

`ifndef complex_dsp

//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////
// Definition of a 16-bit floating point multiplier
// This is a heavily modified version of:
// https://github.com/fbrosser/DSP48E1-FP/tree/master/src/FPMult
// Original author: Fredrik Brosser
// Abridged by: Samidh Mehta
//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////

module FPMult_16_systolic_4x4_fp(
		clk,
		rst,
		a,
		b,
		result,
		flags
    );
	
	// Input Ports
	input clk ;							// Clock
	input rst ;							// Reset signal
	input [`DWIDTH-1:0] a;						// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b;						// Input B, a 32-bit floating point number
	
	// Output ports
	output [`DWIDTH-1:0] result ;					// Product, result of the operation, 32-bit FP number
	output [4:0] flags ;						// Flags indicating exceptions according to IEEE754
	
	// Internal signals
	wire [`DWIDTH-1:0] Z_int ;					// Product, result of the operation, 32-bit FP number
	wire [4:0] Flags_int ;						// Flags indicating exceptions according to IEEE754
	
	wire Sa ;							// A's sign
	wire Sb ;							// B's sign
	wire Sp ;							// Product sign
	wire [`EXPONENT-1:0] Ea ;					// A's exponent
	wire [`EXPONENT-1:0] Eb ;					// B's exponent
	wire [2*`MANTISSA+1:0] Mp ;					// Product mantissa
	wire [4:0] InputExc ;						// Exceptions in inputs
	wire [`MANTISSA-1:0] NormM ;					// Normalized mantissa
	wire [`EXPONENT:0] NormE ;					// Normalized exponent
	wire [`MANTISSA:0] RoundM ;					// Normalized mantissa
	wire [`EXPONENT:0] RoundE ;					// Normalized exponent
	wire [`MANTISSA:0] RoundMP ;					// Normalized mantissa
	wire [`EXPONENT:0] RoundEP ;					// Normalized exponent
	wire GRS ;

	//reg [63:0] pipe_0;						// Pipeline register Input->Prep
	reg [2*`DWIDTH-1:0] pipe_0;					// Pipeline register Input->Prep

	//reg [92:0] pipe_1;						// Pipeline register Prep->Execute
	//reg [3*`MANTISSA+2*`EXPONENT+7:0] pipe_1;			// Pipeline register Prep->Execute
	reg [3*`MANTISSA+2*`EXPONENT+18:0] pipe_1;

	//reg [38:0] pipe_2;						// Pipeline register Execute->Normalize
	reg [`MANTISSA+`EXPONENT+7:0] pipe_2;				// Pipeline register Execute->Normalize
	
	//reg [72:0] pipe_3;						// Pipeline register Normalize->Round
	reg [2*`MANTISSA+2*`EXPONENT+10:0] pipe_3;			// Pipeline register Normalize->Round

	//reg [36:0] pipe_4;						// Pipeline register Round->Output
	reg [`DWIDTH+4:0] pipe_4;					// Pipeline register Round->Output
	
	assign result = pipe_4[`DWIDTH+4:5] ;
	assign flags = pipe_4[4:0] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPMult_PrepModule_systolic_4x4_fp PrepModule(clk, rst, pipe_0[2*`DWIDTH-1:`DWIDTH], pipe_0[`DWIDTH-1:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA+1:0], InputExc[4:0]) ;

	// Perform (unsigned) mantissa multiplication
	FPMult_ExecuteModule_systolic_4x4_fp ExecuteModule(pipe_1[3*`MANTISSA+`EXPONENT*2+7:2*`MANTISSA+2*`EXPONENT+8], pipe_1[2*`MANTISSA+2*`EXPONENT+7:2*`MANTISSA+7], pipe_1[2*`MANTISSA+6:5], pipe_1[2*`MANTISSA+2*`EXPONENT+6:2*`MANTISSA+`EXPONENT+7], pipe_1[2*`MANTISSA+`EXPONENT+6:2*`MANTISSA+7], pipe_1[2*`MANTISSA+2*`EXPONENT+8], pipe_1[2*`MANTISSA+2*`EXPONENT+7], Sp, NormE[`EXPONENT:0], NormM[`MANTISSA-1:0], GRS) ;

	// Round result and if necessary, perform a second (post-rounding) normalization step
	FPMult_NormalizeModule_systolic_4x4_fp NormalizeModule(pipe_2[`MANTISSA-1:0], pipe_2[`MANTISSA+`EXPONENT:`MANTISSA], RoundE[`EXPONENT:0], RoundEP[`EXPONENT:0], RoundM[`MANTISSA:0], RoundMP[`MANTISSA:0]) ;		

	// Round result and if necessary, perform a second (post-rounding) normalization step
	//FPMult_RoundModule_systolic_4x4_fp RoundModule(pipe_3[47:24], pipe_3[23:0], pipe_3[65:57], pipe_3[56:48], pipe_3[66], pipe_3[67], pipe_3[72:68], Z_int[31:0], Flags_int[4:0]) ;		
	FPMult_RoundModule_systolic_4x4_fp RoundModule(pipe_3[2*`MANTISSA+1:`MANTISSA+1], pipe_3[`MANTISSA:0], pipe_3[2*`MANTISSA+2*`EXPONENT+3:2*`MANTISSA+`EXPONENT+3], pipe_3[2*`MANTISSA+`EXPONENT+2:2*`MANTISSA+2], pipe_3[2*`MANTISSA+2*`EXPONENT+4], pipe_3[2*`MANTISSA+2*`EXPONENT+5], pipe_3[2*`MANTISSA+2*`EXPONENT+10:2*`MANTISSA+2*`EXPONENT+6], Z_int[`DWIDTH-1:0], Flags_int[4:0]) ;		

//adding always@ (*) instead of posedge clock to make design combinational
	always @ (posedge clk) begin	
		if(rst) begin
			pipe_0 <= 0;
			pipe_1 <= 0;
			pipe_2 <= 0; 
			pipe_3 <= 0;
			pipe_4 <= 0;
		end 
		else begin		
			/* PIPE 0
				[2*`DWIDTH-1:`DWIDTH] A
				[`DWIDTH-1:0] B
			*/
                       pipe_0 <= {a, b} ;


			/* PIPE 1
				[2*`EXPONENT+3*`MANTISSA + 18: 2*`EXPONENT+2*`MANTISSA + 18] //pipe_0[`DWIDTH+`MANTISSA-1:`DWIDTH] , mantissa of A
				[2*`EXPONENT+2*`MANTISSA + 17 :2*`EXPONENT+2*`MANTISSA + 9] // pipe_0[8:0]
				[2*`EXPONENT+2*`MANTISSA + 8] Sa
				[2*`EXPONENT+2*`MANTISSA + 7] Sb
				[2*`EXPONENT+2*`MANTISSA + 6:`EXPONENT+2*`MANTISSA+7] Ea
				[`EXPONENT +2*`MANTISSA+6:2*`MANTISSA+7] Eb
				[2*`MANTISSA+1+5:5] Mp
				[4:0] InputExc
			*/
			//pipe_1 <= {pipe_0[`DWIDTH+`MANTISSA-1:`DWIDTH], pipe_0[`MANTISSA_MUL_SPLIT_LSB-1:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA-1:0], InputExc[4:0]} ;
			pipe_1 <= {pipe_0[`DWIDTH+`MANTISSA-1:`DWIDTH], pipe_0[8:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA+1:0], InputExc[4:0]} ;
			
			/* PIPE 2
				[`EXPONENT + `MANTISSA + 7:`EXPONENT + `MANTISSA + 3] InputExc
				[`EXPONENT + `MANTISSA + 2] GRS
				[`EXPONENT + `MANTISSA + 1] Sp
				[`EXPONENT + `MANTISSA:`MANTISSA] NormE
				[`MANTISSA-1:0] NormM
			*/
			pipe_2 <= {pipe_1[4:0], GRS, Sp, NormE[`EXPONENT:0], NormM[`MANTISSA-1:0]} ;
			/* PIPE 3
				[2*`EXPONENT+2*`MANTISSA+10:2*`EXPONENT+2*`MANTISSA+6] InputExc
				[2*`EXPONENT+2*`MANTISSA+5] GRS
				[2*`EXPONENT+2*`MANTISSA+4] Sp	
				[2*`EXPONENT+2*`MANTISSA+3:`EXPONENT+2*`MANTISSA+3] RoundE
				[`EXPONENT+2*`MANTISSA+2:2*`MANTISSA+2] RoundEP
				[2*`MANTISSA+1:`MANTISSA+1] RoundM
				[`MANTISSA:0] RoundMP
			*/
			pipe_3 <= {pipe_2[`EXPONENT+`MANTISSA+7:`EXPONENT+`MANTISSA+1], RoundE[`EXPONENT:0], RoundEP[`EXPONENT:0], RoundM[`MANTISSA:0], RoundMP[`MANTISSA:0]} ;
			/* PIPE 4
				[`DWIDTH+4:5] Z
				[4:0] Flags
			*/				
			pipe_4 <= {Z_int[`DWIDTH-1:0], Flags_int[4:0]} ;
		end
	end
		
endmodule



module FPMult_PrepModule_systolic_4x4_fp (
		clk,
		rst,
		a,
		b,
		Sa,
		Sb,
		Ea,
		Eb,
		Mp,
		InputExc
	);
	
	// Input ports
	input clk ;
	input rst ;
	input [`DWIDTH-1:0] a ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b ;								// Input B, a 32-bit floating point number
	
	// Output ports
	output Sa ;										// A's sign
	output Sb ;										// B's sign
	output [`EXPONENT-1:0] Ea ;								// A's exponent
	output [`EXPONENT-1:0] Eb ;								// B's exponent
	output [2*`MANTISSA+1:0] Mp ;							// Mantissa product
	output [4:0] InputExc ;						// Input numbers are exceptions
	
	// Internal signals							// If signal is high...
	wire ANaN ;										// A is a signalling NaN
	wire BNaN ;										// B is a signalling NaN
	wire AInf ;										// A is infinity
	wire BInf ;										// B is infinity
    wire [`MANTISSA-1:0] Ma;
    wire [`MANTISSA-1:0] Mb;
	
	assign ANaN = &(a[`DWIDTH-2:`MANTISSA]) &  |(a[`DWIDTH-2:`MANTISSA]) ;			// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(b[`DWIDTH-2:`MANTISSA]) &  |(b[`MANTISSA-1:0]);			// All one exponent and not all zero mantissa - NaN
	assign AInf = &(a[`DWIDTH-2:`MANTISSA]) & ~|(a[`DWIDTH-2:`MANTISSA]) ;		// All one exponent and all zero mantissa - Infinity
	assign BInf = &(b[`DWIDTH-2:`MANTISSA]) & ~|(b[`DWIDTH-2:`MANTISSA]) ;		// All one exponent and all zero mantissa - Infinity
	
	// Check for any exceptions and put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	//assign InputExc = {(ANaN | ANaN | BNaN |BNaN), ANaN, ANaN, BNaN,BNaN} ;
	
	// Take input numbers apart
	assign Sa = a[`DWIDTH-1] ;							// A's sign
	assign Sb = b[`DWIDTH-1] ;							// B's sign
	assign Ea = a[`DWIDTH-2:`MANTISSA];						// Store A's exponent in Ea, unless A is an exception
	assign Eb = b[`DWIDTH-2:`MANTISSA];						// Store B's exponent in Eb, unless B is an exception	
//    assign Ma = a[`MANTISSA_MSB:`MANTISSA_LSB];
  //  assign Mb = b[`MANTISSA_MSB:`MANTISSA_LSB];
	


	//assign Mp = ({4'b0001, a[`MANTISSA-1:0]}*{4'b0001, b[`MANTISSA-1:9]}) ;
	assign Mp = ({1'b1,a[`MANTISSA-1:0]}*{1'b1, b[`MANTISSA-1:0]}) ;

	
    //We multiply part of the mantissa here
    //Full mantissa of A
    //Bits MANTISSA_MUL_SPLIT_MSB:MANTISSA_MUL_SPLIT_LSB of B
   // wire [`ACTUAL_MANTISSA-1:0] inp_A;
   // wire [`ACTUAL_MANTISSA-1:0] inp_B;
   // assign inp_A = {1'b1, Ma};
   // assign inp_B = {{(`MANTISSA-(`MANTISSA_MUL_SPLIT_MSB-`MANTISSA_MUL_SPLIT_LSB+1)){1'b0}}, 1'b1, Mb[`MANTISSA_MUL_SPLIT_MSB:`MANTISSA_MUL_SPLIT_LSB]};
   // DW02_mult #(`ACTUAL_MANTISSA,`ACTUAL_MANTISSA) u_mult(.A(inp_A), .B(inp_B), .TC(1'b0), .PRODUCT(Mp));
endmodule


module FPMult_ExecuteModule_systolic_4x4_fp(
		a,
		b,
		MpC,
		Ea,
		Eb,
		Sa,
		Sb,
		Sp,
		NormE,
		NormM,
		GRS
    );

	// Input ports
	input [`MANTISSA-1:0] a ;
	input [2*`EXPONENT:0] b ;
	input [2*`MANTISSA+1:0] MpC ;
	input [`EXPONENT-1:0] Ea ;						// A's exponent
	input [`EXPONENT-1:0] Eb ;						// B's exponent
	input Sa ;								// A's sign
	input Sb ;								// B's sign
	
	// Output ports
	output Sp ;								// Product sign
	output [`EXPONENT:0] NormE ;													// Normalized exponent
	output [`MANTISSA-1:0] NormM ;												// Normalized mantissa
	output GRS ;
	
	wire [2*`MANTISSA+1:0] Mp ;
	
	assign Sp = (Sa ^ Sb) ;												// Equal signs give a positive product
	
   // wire [`ACTUAL_MANTISSA-1:0] inp_a;
   // wire [`ACTUAL_MANTISSA-1:0] inp_b;
   // assign inp_a = {1'b1, a};
   // assign inp_b = {{(`MANTISSA-`MANTISSA_MUL_SPLIT_LSB){1'b0}}, 1'b0, b};
   // DW02_mult #(`ACTUAL_MANTISSA,`ACTUAL_MANTISSA) u_mult(.A(inp_a), .B(inp_b), .TC(1'b0), .PRODUCT(Mp_temp));
   // DW01_add #(2*`ACTUAL_MANTISSA) u_add(.A(Mp_temp), .B(MpC<<`MANTISSA_MUL_SPLIT_LSB), .CI(1'b0), .SUM(Mp), .CO());

	//assign Mp = (MpC<<(2*`EXPONENT+1)) + ({4'b0001, a[`MANTISSA-1:0]}*{1'b0, b[2*`EXPONENT:0]}) ;
	assign Mp = MpC;


	assign NormM = (Mp[2*`MANTISSA+1] ? Mp[2*`MANTISSA:`MANTISSA+1] : Mp[2*`MANTISSA-1:`MANTISSA]); 	// Check for overflow
	assign NormE = (Ea + Eb + Mp[2*`MANTISSA+1]);								// If so, increment exponent
	
	assign GRS = ((Mp[`MANTISSA]&(Mp[`MANTISSA+1]))|(|Mp[`MANTISSA-1:0])) ;
	
endmodule

module FPMult_NormalizeModule_systolic_4x4_fp(
		NormM,
		NormE,
		RoundE,
		RoundEP,
		RoundM,
		RoundMP
    );

	// Input Ports
	input [`MANTISSA-1:0] NormM ;									// Normalized mantissa
	input [`EXPONENT:0] NormE ;									// Normalized exponent

	// Output Ports
	output [`EXPONENT:0] RoundE ;
	output [`EXPONENT:0] RoundEP ;
	output [`MANTISSA:0] RoundM ;
	output [`MANTISSA:0] RoundMP ; 
	
// EXPONENT = 5 
// EXPONENT -1 = 4
// NEED to subtract 2^4 -1 = 15

wire [`EXPONENT-1 : 0] bias;

assign bias =  ((1<< (`EXPONENT -1)) -1);

	assign RoundE = NormE - bias ;
	assign RoundEP = NormE - bias -1 ;
	assign RoundM = NormM ;
	assign RoundMP = NormM ;

endmodule

module FPMult_RoundModule_systolic_4x4_fp(
		RoundM,
		RoundMP,
		RoundE,
		RoundEP,
		Sp,
		GRS,
		InputExc,
		Z,
		Flags
    );

	// Input Ports
	input [`MANTISSA:0] RoundM ;									// Normalized mantissa
	input [`MANTISSA:0] RoundMP ;									// Normalized exponent
	input [`EXPONENT:0] RoundE ;									// Normalized mantissa + 1
	input [`EXPONENT:0] RoundEP ;									// Normalized exponent + 1
	input Sp ;												// Product sign
	input GRS ;
	input [4:0] InputExc ;
	
	// Output Ports
	output [`DWIDTH-1:0] Z ;										// Final product
	output [4:0] Flags ;
	
	// Internal Signals
	wire [`EXPONENT:0] FinalE ;									// Rounded exponent
	wire [`MANTISSA:0] FinalM;
	wire [`MANTISSA:0] PreShiftM;
	
	assign PreShiftM = GRS ? RoundMP : RoundM ;	// Round up if R and (G or S)
	
	// Post rounding normalization (potential one bit shift> use shifted mantissa if there is overflow)
	assign FinalM = (PreShiftM[`MANTISSA] ? {1'b0, PreShiftM[`MANTISSA:1]} : PreShiftM[`MANTISSA:0]) ;
	
	assign FinalE = (PreShiftM[`MANTISSA] ? RoundEP : RoundE) ; // Increment exponent if a shift was done
	
	assign Z = {Sp, FinalE[`EXPONENT-1:0], FinalM[`MANTISSA-1:0]} ;   // Putting the pieces together
	assign Flags = InputExc[4:0];

endmodule

`endif

 
//////////////////////////////////////////////////////////////////////////
// A floating point 16-bit to floating point 32-bit converter
//////////////////////////////////////////////////////////////////////////
`ifndef complex_dsp
module fp16_to_fp32_systolic_4x4_fp (input [15:0] a , output [31:0] b);

reg [31:0]b_temp;
reg [3:0] j;
reg [3:0] k;
reg [3:0] k_temp;
always @ (*) begin

if ( a [14: 0] == 15'b0 ) begin //signed zero
	b_temp [31] = a[15]; //sign bit
	b_temp[30:0] = 31'b0;
end

else begin

	if ( a[14 : 10] == 5'b0 ) begin //denormalized (covert to normalized)
		
		for (j=0; j<=9; j=j+1) begin
			if (a[j] == 1'b1) begin 
			    k_temp = j;	
			end
		end
	k = 9 - k_temp;

	b_temp [22:0] = ( (a [9:0] << (k+1'b1)) & 10'h3FF ) << 13;
	b_temp [30:23] =  7'd127 - 4'd15 - k;
	b_temp [31] = a[15];
	end

	else if ( a[14 : 10] == 5'b11111 ) begin //Infinity/ NAN
	b_temp [22:0] = a [9:0] << 13;
	b_temp [30:23] = 8'hFF;
	b_temp [31] = a[15];
	end

	else begin //Normalized Number
	b_temp [22:0] = a [9:0] << 13;
	b_temp [30:23] =  7'd127 - 4'd15 + a[14:10];
	b_temp [31] = a[15];
	end
end
end

assign b = b_temp;


endmodule

//////////////////////////////////////////////////////////////////////////
// A floating point 32-bit to floating point 16-bit converter
//////////////////////////////////////////////////////////////////////////
module fp32_to_fp16_systolic_4x4_fp (input [31:0] a , output [15:0] b);

reg [15:0]b_temp;
//integer j;
//reg [3:0]k;
always @ (*) begin

if ( a [30: 0] == 15'b0 ) begin //signed zero
	b_temp [15] = a[30]; //sign bit
	b_temp [14:0] = 15'b0; 
end

else begin

	if ( a[30 : 23] <= 8'd112  &&  a[30 : 23] >= 8'd103 ) begin //denormalized (covert to normalized)
		
	b_temp [9:0] = {1'b1, a[22:13]} >> {8'd112 - a[30 : 23] + 1'b1} ;  
	b_temp [14:10] =  5'b0;
	b_temp [15] = a[31];
	end

	else if ( a[ 30 : 23] == 8'b11111111 ) begin //Infinity/ NAN
	b_temp [9:0] = a [22:13];
	b_temp [14:10] = 5'h1F;
	b_temp [15] = a[31];
	end

	else begin //Normalized Number
	b_temp [9:0] = a [22:13];
	b_temp [14:10] = 4'd15 - 7'd127  + a[30:23]; //number should be in the range which can be depicted by fp16 (exp for fp32: 70h, 8Eh ; normalized exp for fp32: -15 to 15)
	b_temp [15] = a[31];
	end
end
end

assign b = b_temp;


endmodule
`endif

//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////
// Definition of a 32-bit floating point adder/subtractor
// This is a heavily modified version of:
// https://github.com/fbrosser/DSP48E1-FP/tree/master/src/FP_AddSub
// Original author: Fredrik Brosser
// Abridged by: Samidh Mehta
//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////

`ifndef complex_dsp
module FPAddSub_single_systolic_4x4_fp(
		clk,
		rst,
		a,
		b,
		operation,
		result,
		flags
	);

// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [31:0] a ;								// Input A, a 32-bit floating point number
	input [31:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [31:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754

	reg [68:0]pipe_1;
	reg [54:0]pipe_2;
	reg [45:0]pipe_3;


//internal module wires

//output ports
	wire Opout;
	wire Sa;
	wire Sb;
	wire MaxAB;
	wire [7:0] CExp;
	wire [4:0] Shift;
	wire [22:0] Mmax;
	wire [4:0] InputExc;
	wire [23:0] Mmin_3;

	wire [32:0] SumS_5 ;
	wire [4:0] Shift_1;							
	wire PSgn ;							
	wire Opr ;	
	
	wire [22:0] NormM ;				// Normalized mantissa
	wire [8:0] NormE ;					// Adjusted exponent
	wire ZeroSum ;						// Zero flag
	wire NegE ;							// Flag indicating negative exponent
	wire R ;								// Round bit
	wire S ;								// Final sticky bit
	wire FG ;

FPAddSub_a_systolic_4x4_fp M1(a,b,operation,Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3);

FPAddSub_b_systolic_4x4_fp M2(pipe_1[51:29],pipe_1[23:0],pipe_1[67],pipe_1[66],pipe_1[65],pipe_1[68],SumS_5,Shift_1,PSgn,Opr);

FPAddSub_c_systolic_4x4_fp M3(pipe_2[54:22],pipe_2[21:17],pipe_2[16:9],NormM,NormE,ZeroSum,NegE,R,S,FG);

FPAddSub_d_systolic_4x4_fp M4(pipe_3[13],pipe_3[22:14],pipe_3[45:23],pipe_3[11],pipe_3[10],pipe_3[9],pipe_3[8],pipe_3[7],pipe_3[6],pipe_3[5],pipe_3[12],pipe_3[4:0],result,flags );


always @ (posedge clk) begin	
		if(rst) begin
			pipe_1 <= 0;
			pipe_2 <= 0;
			pipe_3 <= 0;
		end 
		else begin
/*
pipe_1:
	[68] Opout;
	[67] Sa;
	[66] Sb;
	[65] MaxAB;
	[64:57] CExp;
	[56:52] Shift;
	[51:29] Mmax;
	[28:24] InputExc;
	[23:0] Mmin_3;	
*/

pipe_1 <= {Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3};

/*
pipe_2:
	[54:22]SumS_5;
	[21:17]Shift;
	[16:9]CExp;	
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_2 <= {SumS_5,Shift_1,pipe_1[64:57], pipe_1[67], pipe_1[66], pipe_1[68], pipe_1[65], pipe_1[28:24] };

/*
pipe_3:
	[45:23] NormM ;				
	[22:14] NormE ;					
	[13]ZeroSum ;						
	[12]NegE ;							
	[11]R ;								
	[10]S ;								
	[9]FG ;
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_3 <= {NormM,NormE,ZeroSum,NegE,R,S,FG, pipe_2[8], pipe_2[7], pipe_2[6], pipe_2[5], pipe_2[4:0] };

end
end

endmodule

// Prealign + Align + Shift 1 + Shift 2
module FPAddSub_a_systolic_4x4_fp(
		A,
		B,
		operation,
		Opout,
		Sa,
		Sb,
		MaxAB,
		CExp,
		Shift,
		Mmax,
		InputExc,
		Mmin_3
		
		
	);
	
	// Input ports
	input [31:0] A ;										// Input A, a 32-bit floating point number
	input [31:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	//output ports
	output Opout;
	output Sa;
	output Sb;
	output MaxAB;
	output [7:0] CExp;
	output [4:0] Shift;
	output [22:0] Mmax;
	output [4:0] InputExc;
	output [23:0] Mmin_3;	
							
	wire [9:0] ShiftDet ;							
	wire [30:0] Aout ;
	wire [30:0] Bout ;
	

	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [7:0] DAB ;										// ExpA - ExpB					
	wire [7:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[30:23]) & |(A[22:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[30:23]) & |(B[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[30:23]) & ~|(A[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[30:23]) & ~|(B[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
  assign DAB = (A[30:23] + ~(B[30:23]) + 1) ;
	assign DBA = (B[30:23] + ~(A[30:23]) + 1) ;

	assign Sa = A[31] ;									// A's sign bit
	assign Sb = B[31] ;									// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[30:0] ;
	assign Bout = B[30:0] ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Output ports
													// Number of steps to smaller mantissa shift right
	wire [22:0] Mmin_1 ;							// Smaller mantissa 
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (Aout[30:0] < Bout[30:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[9:5] : ShiftDet[4:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin_1 = MaxAB ? Aout[22:0] : Bout[22:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? Bout[22:0]: Aout[22:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? Bout[30:23] : Aout[30:23]) ;	

// Input ports
					// Smaller mantissa after 16|12|8|4 shift
	wire [2:0] Shift_1 ;						// Shift amount
	
	assign Shift_1 = Shift [4:2];

	wire [23:0] Mmin_2 ;						// The smaller mantissa
	
	// Internal signals
	reg	  [23:0]		Lvl1;
	reg	  [23:0]		Lvl2;
	wire    [47:0]    Stage1;	
	integer           i;                // Loop variable
	
	always @(*) begin						
		// Rotate by 16?
		Lvl1 <= Shift_1[2] ? {17'b00000000000000001, Mmin_1[22:16]} : {1'b1, Mmin_1}; 
	end
	
	assign Stage1 = {Lvl1, Lvl1};
	
	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift_1[1:0])
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[23:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[23:19] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[23:15] <= 0; end
			// Rotate by 12	
			2'b11:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[23:11] <= 0; end
	  endcase
	end
	
	// Assign output to next shift stage
	assign Mmin_2 = Lvl2;
								// Smaller mantissa after 16|12|8|4 shift
	wire [1:0] Shift_2 ;						// Shift amount
	
	assign Shift_2 =Shift  [1:0] ;
					// The smaller mantissa
	
	// Internal Signal
	reg	  [23:0]		Lvl3;
	wire    [47:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {Mmin_2, Mmin_2};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_2[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[23:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[23] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[23:22] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[23:21] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin_3 = Lvl3;	

	
endmodule

module FPAddSub_b_systolic_4x4_fp(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		SumS_5,
		Shift,
		PSgn,
		Opr
);
	input [22:0] Mmax ;					// The larger mantissa
	input [23:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	wire [32:0] Sum ;	
						// Output ports
	output [32:0] SumS_5 ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount				// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation

	// Perform effective operation
	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, 8'b00000000} - {Mmin, 8'b00000000}) : ({1'b1, Mmax, 8'b00000000} + {Mmin, 8'b00000000}) ;
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

		// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[32] ? 5'b00000 :	 
		Sum[31] ? 5'b00001 : 
		Sum[30] ? 5'b00010 : 
		Sum[29] ? 5'b00011 : 
		Sum[28] ? 5'b00100 : 
		Sum[27] ? 5'b00101 : 
		Sum[26] ? 5'b00110 : 
		Sum[25] ? 5'b00111 :
		Sum[24] ? 5'b01000 :
		Sum[23] ? 5'b01001 :
		Sum[22] ? 5'b01010 :
		Sum[21] ? 5'b01011 :
		Sum[20] ? 5'b01100 :
		Sum[19] ? 5'b01101 :
		Sum[18] ? 5'b01110 :
		Sum[17] ? 5'b01111 :
		Sum[16] ? 5'b10000 :
		Sum[15] ? 5'b10001 :
		Sum[14] ? 5'b10010 :
		Sum[13] ? 5'b10011 :
		Sum[12] ? 5'b10100 :
		Sum[11] ? 5'b10101 :
		Sum[10] ? 5'b10110 :
		Sum[9] ? 5'b10111 :
		Sum[8] ? 5'b11000 :
		Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [32:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[16:0], 16'b0000000000000000} : Sum; 
	end
	
	// Assign outputs
	assign SumS_5 = Lvl1;	

endmodule

module FPAddSub_c_systolic_4x4_fp(
		SumS_5,
		Shift,
		CExp,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [32:0] SumS_5 ;						// Smaller mantissa after 16|12|8|4 shift
	
	input [4:0] Shift ;						// Shift amount
	
// Input ports
	
	input [7:0] CExp ;
	

	// Output ports
	output [22:0] NormM ;				// Normalized mantissa
	output [8:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;


	wire [3:0]Shift_1;
	assign Shift_1 = Shift [3:0];
	// Output ports
	wire [32:0] SumS_7 ;						// The smaller mantissa
	
	reg	  [32:0]		Lvl2;
	wire    [65:0]    Stage1;	
	reg	  [32:0]		Lvl3;
	wire    [65:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {SumS_5, SumS_5};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[32:0];       		
			// Rotate by 4
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_1[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[32:0];
			// Rotate by 1
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign SumS_7 = Lvl3;						// Take out smaller mantissa



	
	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [8:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [8:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = SumS_7[32] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|SumS_7 ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[8] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = SumS_7[31:9] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = SumS_7[8] ; 
	assign R = SumS_7[7] ;
	assign S = |SumS_7[6:0] ;		
	
endmodule

module FPAddSub_d_systolic_4x4_fp(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		NegE,
		InputExc,
		P,
		Flags 
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [8:0] NormE ;				// Normalized exponent
	input [22:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	

	input NegE ;						// Negative exponent?
	input [4:0] InputExc ;					// Exceptions in inputs A and B

	// Output ports
	output [31:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// 
	wire [31:0] Z ;					// Final result
	wire EOF ;
	
	// Internal signals
	wire [23:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [22:0] RoundM ;				// The final rounded sum
	wire [8:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	wire FSgn;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[22:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[23] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? 8'b00000000 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[7:0], RoundM[22:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[8];

/////////////////////////////////////////////////////////////////////////////////////////////////////////



	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[30:23]) & ~|(Z[30:23]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule
`endif

module spram_4096_60bit (
    clk,
    address,
    wren,
    data,
    out
);
parameter AWIDTH=12;
parameter NUM_WORDS=4096;
parameter DWIDTH=60;
input clk;
input [(AWIDTH-1):0] address;
input  wren;
input [(DWIDTH-1):0] data;
output reg [(DWIDTH-1):0] out;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren) begin
      ram[address] <= data;
  end
  else begin
      out <= ram[address];
  end
end
  
`else

defparam u_single_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_single_port_ram.DATA_WIDTH = DWIDTH;

single_port_ram u_single_port_ram(
.addr(address),
.we(wren),
.data(data),
.out(out),
.clk(clk)
);

`endif

endmodule

module adder_tree_4stage_8bit(clk,reset,inp00,inp01,inp10,inp11,inp20,inp21,inp30,inp31,inp40,inp41,inp50,inp51,inp60,inp61,inp70,inp71,sum_out);

input clk;
input reset; 
input [7:0] inp00; 
input [7:0] inp01;
input [7:0] inp10; 
input [7:0] inp11;
input [7:0] inp20; 
input [7:0] inp21;
input [7:0] inp30; 
input [7:0] inp31;
input [7:0] inp40; 
input [7:0] inp41;
input [7:0] inp50; 
input [7:0] inp51;
input [7:0] inp60; 
input [7:0] inp61;
input [7:0] inp70; 
input [7:0] inp71;
output reg [15:0] sum_out;

reg [8:0] S_0_0; 
reg [8:0] S_0_1;
reg [8:0] S_0_2;
reg [8:0] S_0_3;
reg [8:0] S_0_4;
reg [8:0] S_0_5;
reg [8:0] S_0_6;
reg [8:0] S_0_7;

always@(posedge clk) begin 

S_0_0 <= inp00 + inp01; 
S_0_1 <= inp10 + inp11;
S_0_2 <= inp20 + inp21;
S_0_3 <= inp30 + inp31;
S_0_4 <= inp40 + inp41; 
S_0_5 <= inp50 + inp51;
S_0_6 <= inp60 + inp61;
S_0_7 <= inp70 + inp71;

end 

reg [9:0] S_1_0;
reg [9:0] S_1_1;
reg [9:0] S_1_2;
reg [9:0] S_1_3;

always@(posedge clk) begin 

S_1_0 <= S_0_0 + S_0_1; 
S_1_1 <= S_0_2 + S_0_3;
S_1_2 <= S_0_4 + S_0_5; 
S_1_3 <= S_0_6 + S_0_7;

end

reg [10:0] S_2_0; 
reg [10:0] S_2_1;

always@(posedge clk) begin 

S_2_0 <= S_1_0 + S_1_1; 
S_2_1 <= S_1_2 + S_1_3;

end

always@(posedge clk) begin 

if (reset == 1'b1) begin 
  sum_out <= 16'd0; 
end
else begin 
  sum_out <= S_2_0 + S_2_1; 
end

end 

endmodule
module spram_4096_40bit (
    clk,
    address,
    wren,
    data,
    out
);
parameter AWIDTH=12;
parameter NUM_WORDS=4096;
parameter DWIDTH=40;
input clk;
input [(AWIDTH-1):0] address;
input  wren;
input [(DWIDTH-1):0] data;
output reg [(DWIDTH-1):0] out;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren) begin
      ram[address] <= data;
  end
  else begin
      out <= ram[address];
  end
end
  
`else

defparam u_single_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_single_port_ram.DATA_WIDTH = DWIDTH;

single_port_ram u_single_port_ram(
.addr(address),
.we(wren),
.data(data),
.out(out),
.clk(clk)
);

`endif

endmodule

`define EXPONENT 5
`define MANTISSA 10
`define ACTUAL_MANTISSA 11
`define EXPONENT_LSB 10
`define EXPONENT_MSB 14
`define MANTISSA_LSB 0
`define MANTISSA_MSB 9
`define MANTISSA_MUL_SPLIT_LSB 3
`define MANTISSA_MUL_SPLIT_MSB 9
`define SIGN 1
`define SIGN_LOC 15
`define DWIDTH (`SIGN+`EXPONENT+`MANTISSA)
`define IEEE_COMPLIANCE 1
`define DATAWIDTH 16

module mode4_adder_tree(
  inp0, 
  inp1, 
  inp2, 
  inp3, 
  inp4, 
  inp5, 
  inp6, 
  inp7, 
  mode4_stage0_run,
  mode4_stage1_run,
  mode4_stage2_run,
  mode4_stage3_run,

  clk,
  reset,
  outp
);

  input clk;
  input reset;
  input  [`DATAWIDTH-1 : 0] inp0; 
  input  [`DATAWIDTH-1 : 0] inp1; 
  input  [`DATAWIDTH-1 : 0] inp2; 
  input  [`DATAWIDTH-1 : 0] inp3; 
  input  [`DATAWIDTH-1 : 0] inp4; 
  input  [`DATAWIDTH-1 : 0] inp5; 
  input  [`DATAWIDTH-1 : 0] inp6; 
  input  [`DATAWIDTH-1 : 0] inp7; 
  output [`DATAWIDTH-1 : 0] outp;
  input mode4_stage0_run;
  input mode4_stage1_run;
  input mode4_stage2_run;
  input mode4_stage3_run;

  wire   [`DATAWIDTH-1 : 0] add0_out_stage3;
  reg    [`DATAWIDTH-1 : 0] add0_out_stage3_reg;
  wire   [`DATAWIDTH-1 : 0] add1_out_stage3;
  reg    [`DATAWIDTH-1 : 0] add1_out_stage3_reg;
  wire   [`DATAWIDTH-1 : 0] add2_out_stage3;
  reg    [`DATAWIDTH-1 : 0] add2_out_stage3_reg;
  wire   [`DATAWIDTH-1 : 0] add3_out_stage3;
  reg    [`DATAWIDTH-1 : 0] add3_out_stage3_reg;

  wire   [`DATAWIDTH-1 : 0] add0_out_stage2;
  reg    [`DATAWIDTH-1 : 0] add0_out_stage2_reg;
  wire   [`DATAWIDTH-1 : 0] add1_out_stage2;
  reg    [`DATAWIDTH-1 : 0] add1_out_stage2_reg;

  wire   [`DATAWIDTH-1 : 0] add0_out_stage1;
  reg    [`DATAWIDTH-1 : 0] add0_out_stage1_reg;

  wire   [`DATAWIDTH-1 : 0] add0_out_stage0;
  reg    [`DATAWIDTH-1 : 0] outp;

//  always @(posedge clk) begin
//    if (reset) begin
//      outp <= 0;
//      add0_out_stage3_reg <= 0;
//      add1_out_stage3_reg <= 0;
//      add2_out_stage3_reg <= 0;
//      add3_out_stage3_reg <= 0;
//      add0_out_stage2_reg <= 0;
//      add1_out_stage2_reg <= 0;
//      add0_out_stage1_reg <= 0;
//    end
//
//    if(~reset && mode4_stage3_run) begin
//      add0_out_stage3_reg <= add0_out_stage3;
//      add1_out_stage3_reg <= add1_out_stage3;
//      add2_out_stage3_reg <= add2_out_stage3;
//      add3_out_stage3_reg <= add3_out_stage3;
//    end
//
//    if(~reset && mode4_stage2_run) begin
//      add0_out_stage2_reg <= add0_out_stage2;
//      add1_out_stage2_reg <= add1_out_stage2;
//    end
//
//    if(~reset && mode4_stage1_run) begin
//      add0_out_stage1_reg <= add0_out_stage1;
//    end
//
//    if(~reset && mode4_stage0_run) begin
//      outp <= add0_out_stage0;
//    end
//
//  end


always @ (posedge clk) begin
	if(~reset && mode4_stage3_run) begin
      add0_out_stage3_reg <= add0_out_stage3;
      add1_out_stage3_reg <= add1_out_stage3;
      add2_out_stage3_reg <= add2_out_stage3;
      add3_out_stage3_reg <= add3_out_stage3;
    end
	
	else if (reset) begin
		add0_out_stage3_reg <= 0;
		add1_out_stage3_reg <= 0;
		add2_out_stage3_reg <= 0;
		add3_out_stage3_reg <= 0;
	end
end		

always @ (posedge clk) begin
	if(~reset && mode4_stage2_run) begin
      add0_out_stage2_reg <= add0_out_stage2;
      add1_out_stage2_reg <= add1_out_stage2;
    end
	
	else if (reset) begin
		add0_out_stage2_reg <= 0;
		add1_out_stage2_reg <= 0;
	end
end		

always @ (posedge clk) begin
	if(~reset && mode4_stage1_run) begin
      add0_out_stage1_reg <= add0_out_stage1;
    end
	else if (reset) begin
	add0_out_stage1_reg <= 0;
	end
end

always @ (posedge clk) begin
	if(~reset && mode4_stage0_run) begin
		outp <= add0_out_stage0;
    end
	else if (reset) begin
		outp <= 0;
	end
end	

  wire clk_NC;
  wire rst_NC;
  wire [4:0] flags_NC0, flags_NC1, flags_NC2, flags_NC3;
  wire [4:0] flags_NC4, flags_NC5, flags_NC6, flags_NC7;

  // 0 add, 1 sub
  FPAddSub add0_stage3(.clk(clk), .rst(reset), .a(inp0),	.b(inp1), .operation(1'b0),	.result(add0_out_stage3), .flags(flags_NC0));
  FPAddSub add1_stage3(.clk(clk), .rst(reset), .a(inp2),	.b(inp3), .operation(1'b0),	.result(add1_out_stage3), .flags(flags_NC1));
  FPAddSub add2_stage3(.clk(clk), .rst(reset), .a(inp4),	.b(inp5), .operation(1'b0),	.result(add2_out_stage3), .flags(flags_NC2));
  FPAddSub add3_stage3(.clk(clk), .rst(reset), .a(inp6),	.b(inp7), .operation(1'b0),	.result(add3_out_stage3), .flags(flags_NC3));

  FPAddSub add0_stage2(.clk(clk), .rst(reset), .a(add0_out_stage3_reg),	.b(add1_out_stage3_reg), .operation(1'b0),	.result(add0_out_stage2), .flags(flags_NC4));
  FPAddSub add1_stage2(.clk(clk), .rst(reset), .a(add2_out_stage3_reg),	.b(add3_out_stage3_reg), .operation(1'b0),	.result(add1_out_stage2), .flags(flags_NC5));

  FPAddSub add0_stage1(.clk(clk), .rst(reset), .a(add0_out_stage2_reg),	.b(add1_out_stage2_reg), .operation(1'b0),	.result(add0_out_stage1), .flags(flags_NC6));

  FPAddSub add0_stage0(.clk(clk), .rst(reset), .a(outp),	.b(add0_out_stage1_reg), .operation(1'b0),	.result(add0_out_stage0), .flags(flags_NC7));


//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add0_stage3(.a(inp0),       .b(inp1),      .z(add0_out_stage3), .rnd(3'b000),    .status());
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add1_stage3(.a(inp2),       .b(inp3),      .z(add1_out_stage3), .rnd(3'b000),    .status());
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add2_stage3(.a(inp4),       .b(inp5),      .z(add2_out_stage3), .rnd(3'b000),    .status());
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add3_stage3(.a(inp6),       .b(inp7),      .z(add3_out_stage3), .rnd(3'b000),    .status());
//
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add0_stage2(.a(add0_out_stage3_reg),       .b(add1_out_stage3_reg),      .z(add0_out_stage2), .rnd(3'b000),    .status());
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add1_stage2(.a(add2_out_stage3_reg),       .b(add3_out_stage3_reg),      .z(add1_out_stage2), .rnd(3'b000),    .status());
//
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add0_stage1(.a(add0_out_stage2_reg),       .b(add1_out_stage2_reg),      .z(add0_out_stage1), .rnd(3'b000),    .status());
//
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add0_stage0(.a(outp),       .b(add0_out_stage1_reg),      .z(add0_out_stage0), .rnd(3'b000),    .status());

endmodule

module FPAddSub(
		clk,
		rst,
		a,
		b,
		operation,			// 0 add, 1 sub
		result,
		flags
	);
	
	// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [`DWIDTH-1:0] a ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [`DWIDTH-1:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754
	
	assign flags = 5'b0;
	
//`ifdef complex_dsp
//adder_fp_clk u_add(.clk(clk), .a(a), .b(b),.out(result));
//`else
FPAddSub_16 u_FPAddSub (.clk(clk), .rst(rst), .a(a), .b(b), .operation(1'b0), .result(result), .flags());
//`endif
endmodule

module FPAddSub_16(
		//bf16,
		clk,
		rst,
		a,
		b,
		operation,			// 0 add, 1 sub
		result,
		flags
	);
	//input bf16; //1 for Bfloat16, 0 for IEEE half precision

	// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [`DWIDTH-1:0] a ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [`DWIDTH-1:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754
	
	// Pipeline Registers
	//reg [79:0] pipe_1;							// Pipeline register PreAlign->Align1
	reg [2*`EXPONENT + 2*`DWIDTH + 5:0] pipe_1;							// Pipeline register PreAlign->Align1

	//reg [67:0] pipe_2;							// Pipeline register Align1->Align3
	//reg [2*`EXPONENT+ 2*`MANTISSA + 8:0] pipe_2;							// Pipeline register Align1->Align3
	wire [2*`EXPONENT+ 2*`MANTISSA + 8:0] pipe_2;

	//reg [76:0] pipe_3;	68						// Pipeline register Align1->Align3
	reg [2*`EXPONENT+ 2*`MANTISSA + 9:0] pipe_3;							// Pipeline register Align1->Align3

	//reg [69:0] pipe_4;							// Pipeline register Align3->Execute
	//reg [2*`EXPONENT+ 2*`MANTISSA + 9:0] pipe_4;							// Pipeline register Align3->Execute
	wire [2*`EXPONENT+ 2*`MANTISSA + 9:0] pipe_4;
	
	//reg [51:0] pipe_5;							// Pipeline register Execute->Normalize
	reg [`DWIDTH+`EXPONENT+11:0] pipe_5;							// Pipeline register Execute->Normalize

	//reg [56:0] pipe_6;							// Pipeline register Nomalize->NormalizeShift1
	//reg [`DWIDTH+`EXPONENT+16:0] pipe_6;							// Pipeline register Nomalize->NormalizeShift1
	wire [`DWIDTH+`EXPONENT+16:0] pipe_6;

	//reg [56:0] pipe_7;							// Pipeline register NormalizeShift2->NormalizeShift3
	//reg [`DWIDTH+`EXPONENT+16:0] pipe_7;							// Pipeline register NormalizeShift2->NormalizeShift3
	wire [`DWIDTH+`EXPONENT+16:0] pipe_7;
	//reg [54:0] pipe_8;							// Pipeline register NormalizeShift3->Round
	reg [`EXPONENT*2+`MANTISSA+15:0] pipe_8;							// Pipeline register NormalizeShift3->Round

	//reg [40:0] pipe_9;							// Pipeline register NormalizeShift3->Round
	//reg [`DWIDTH+8:0] pipe_9;							// Pipeline register NormalizeShift3->Round
	wire [`DWIDTH+8:0] pipe_9;

	// Internal wires between modules
	wire [`DWIDTH-2:0] Aout_0 ;							// A - sign
	wire [`DWIDTH-2:0] Bout_0 ;							// B - sign
	wire Opout_0 ;									// A's sign
	wire Sa_0 ;										// A's sign
	wire Sb_0 ;										// B's sign
	wire MaxAB_1 ;									// Indicates the larger of A and B(0/A, 1/B)
	wire [`EXPONENT-1:0] CExp_1 ;							// Common Exponent
	wire [`EXPONENT-1:0] Shift_1 ;							// Number of steps to smaller mantissa shift right (align)
	wire [`MANTISSA-1:0] Mmax_1 ;							// Larger mantissa
	wire [4:0] InputExc_0 ;						// Input numbers are exceptions
	wire [2*`EXPONENT-1:0] ShiftDet_0 ;
	wire [`MANTISSA-1:0] MminS_1 ;						// Smaller mantissa after 0/16 shift
	wire [`MANTISSA:0] MminS_2 ;						// Smaller mantissa after 0/4/8/12 shift
	wire [`MANTISSA:0] Mmin_3 ;							// Smaller mantissa after 0/1/2/3 shift
	wire [`DWIDTH:0] Sum_4 ;
	wire PSgn_4 ;
	wire Opr_4 ;
	wire [`EXPONENT-1:0] Shift_5 ;							// Number of steps to shift sum left (normalize)
	wire [`DWIDTH:0] SumS_5 ;							// Sum after 0/16 shift
	wire [`DWIDTH:0] SumS_6 ;							// Sum after 0/16 shift
	wire [`DWIDTH:0] SumS_7 ;							// Sum after 0/16 shift
	wire [`MANTISSA-1:0] NormM_8 ;						// Normalized mantissa
	wire [`EXPONENT:0] NormE_8;							// Adjusted exponent
	wire ZeroSum_8 ;								// Zero flag
	wire NegE_8 ;									// Flag indicating negative exponent
	wire R_8 ;										// Round bit
	wire S_8 ;										// Final sticky bit
	wire FG_8 ;										// Final sticky bit
	wire [`DWIDTH-1:0] P_int ;
	wire EOF ;
	
	// Prepare the operands for alignment and check for exceptions
	FPAddSub_PrealignModule PrealignModule
	(	// Inputs
		a, b, operation,
		// Outputs
		Sa_0, Sb_0, ShiftDet_0[2*`EXPONENT-1:0], InputExc_0[4:0], Aout_0[`DWIDTH-2:0], Bout_0[`DWIDTH-2:0], Opout_0) ;
		
	// Prepare the operands for alignment and check for exceptions
	FPAddSub_AlignModule AlignModule
	(	// Inputs
		pipe_1[2*`EXPONENT + 2*`DWIDTH + 4: 2*`EXPONENT +`DWIDTH + 6], pipe_1[2*`EXPONENT +`DWIDTH + 5 :  2*`EXPONENT +7], pipe_1[2*`EXPONENT+4:5],
		// Outputs
		CExp_1[`EXPONENT-1:0], MaxAB_1, Shift_1[`EXPONENT-1:0], MminS_1[`MANTISSA-1:0], Mmax_1[`MANTISSA-1:0]) ;	

	// Alignment Shift Stage 1
	FPAddSub_AlignShift1 AlignShift1
	(  // Inputs
		//bf16, 
		pipe_2[`MANTISSA-1:0], pipe_2[`EXPONENT+ 2*`MANTISSA + 4 : 2*`MANTISSA + 7],
		// Outputs
		MminS_2[`MANTISSA:0]) ;

	// Alignment Shift Stage 3 and compution of guard and sticky bits
	FPAddSub_AlignShift2 AlignShift2  
	(  // Inputs
		pipe_3[`MANTISSA:0], pipe_3[2*`MANTISSA+7:2*`MANTISSA+6],
		// Outputs
		Mmin_3[`MANTISSA:0]) ;
						
	// Perform mantissa addition
	FPAddSub_ExecutionModule ExecutionModule
	(  // Inputs
		pipe_4[`MANTISSA*2+5:`MANTISSA+6], pipe_4[`MANTISSA:0], pipe_4[2*`EXPONENT+ 2*`MANTISSA + 8], pipe_4[2*`EXPONENT+ 2*`MANTISSA + 7], pipe_4[2*`EXPONENT+ 2*`MANTISSA + 6], pipe_4[2*`EXPONENT+ 2*`MANTISSA + 9],
		// Outputs
		Sum_4[`DWIDTH:0], PSgn_4, Opr_4) ;
	
	// Prepare normalization of result
	FPAddSub_NormalizeModule NormalizeModule
	(  // Inputs
		pipe_5[`DWIDTH:0], 
		// Outputs
		SumS_5[`DWIDTH:0], Shift_5[4:0]) ;
					
	// Normalization Shift Stage 1
	FPAddSub_NormalizeShift1 NormalizeShift1
	(  // Inputs
		pipe_6[`DWIDTH:0], pipe_6[`DWIDTH+`EXPONENT+14:`DWIDTH+`EXPONENT+11],
		// Outputs
		SumS_7[`DWIDTH:0]) ;
		
	// Normalization Shift Stage 3 and final guard, sticky and round bits
	FPAddSub_NormalizeShift2 NormalizeShift2
	(  // Inputs
		pipe_7[`DWIDTH:0], pipe_7[`DWIDTH+`EXPONENT+5:`DWIDTH+6], pipe_7[`DWIDTH+`EXPONENT+15:`DWIDTH+`EXPONENT+11],
		// Outputs
		NormM_8[`MANTISSA-1:0], NormE_8[`EXPONENT:0], ZeroSum_8, NegE_8, R_8, S_8, FG_8) ;

	// Round and put result together
	FPAddSub_RoundModule RoundModule
	(  // Inputs
		 pipe_8[3], pipe_8[4+`EXPONENT:4], pipe_8[`EXPONENT+`MANTISSA+4:5+`EXPONENT], pipe_8[1], pipe_8[0], pipe_8[`EXPONENT*2+`MANTISSA+15], pipe_8[`EXPONENT*2+`MANTISSA+12], pipe_8[`EXPONENT*2+`MANTISSA+11], pipe_8[`EXPONENT*2+`MANTISSA+14], pipe_8[`EXPONENT*2+`MANTISSA+10], 
		// Outputs
		P_int[`DWIDTH-1:0], EOF) ;
	
	// Check for exceptions
	FPAddSub_ExceptionModule Exceptionmodule
	(  // Inputs
		pipe_9[8+`DWIDTH:9], pipe_9[8], pipe_9[7], pipe_9[6], pipe_9[5:1], pipe_9[0], 
		// Outputs
		result[`DWIDTH-1:0], flags[4:0]) ;			
	

assign pipe_2 = {pipe_1[2*`EXPONENT + 2*`DWIDTH + 5], pipe_1[2*`EXPONENT +6:2*`EXPONENT +5], MaxAB_1, CExp_1[`EXPONENT-1:0], Shift_1[`EXPONENT-1:0], Mmax_1[`MANTISSA-1:0], pipe_1[4:0], MminS_1[`MANTISSA-1:0]} ;
assign pipe_4 = {pipe_3[2*`EXPONENT+ 2*`MANTISSA + 9:`MANTISSA+1], Mmin_3[`MANTISSA:0]} ;
assign pipe_6 = {pipe_5[`DWIDTH+`EXPONENT+11], Shift_5[4:0], pipe_5[`DWIDTH+`EXPONENT+10:`DWIDTH+1], SumS_5[`DWIDTH:0]} ;
assign pipe_7 = {pipe_6[`DWIDTH+`EXPONENT+16:`DWIDTH+1], SumS_7[`DWIDTH:0]} ;
assign pipe_9 = {P_int[`DWIDTH-1:0], pipe_8[2], pipe_8[1], pipe_8[0], pipe_8[`EXPONENT+`MANTISSA+9:`EXPONENT+`MANTISSA+5], EOF} ;

	always @ (posedge clk) begin	
		if(rst) begin
			pipe_1 <= 0;
			//pipe_2 <= 0;
			pipe_3 <= 0;
			//pipe_4 <= 0;
			pipe_5 <= 0;
			//pipe_6 <= 0;
			//pipe_7 <= 0;
			pipe_8 <= 0;
			//pipe_9 <= 0;
		end 
		else begin
/* PIPE_1:
	[2*`EXPONENT + 2*`DWIDTH + 5]  Opout_0
	[2*`EXPONENT + 2*`DWIDTH + 4: 2*`EXPONENT +`DWIDTH + 6] A_out0
	[2*`EXPONENT +`DWIDTH + 5 :  2*`EXPONENT +7] Bout_0
	[2*`EXPONENT +6] Sa_0
	[2*`EXPONENT +5] Sb_0
	[2*`EXPONENT +4 : 5] ShiftDet_0
	[4:0] Input Exc
*/
			pipe_1 <= {Opout_0, Aout_0[`DWIDTH-2:0], Bout_0[`DWIDTH-2:0], Sa_0, Sb_0, ShiftDet_0[2*`EXPONENT -1:0], InputExc_0[4:0]} ;	
/* PIPE_2
[2*`EXPONENT+ 2*`MANTISSA + 8] operation
[2*`EXPONENT+ 2*`MANTISSA + 7] Sa_0
[2*`EXPONENT+ 2*`MANTISSA + 6] Sb_0
[2*`EXPONENT+ 2*`MANTISSA + 5] MaxAB_0
[2*`EXPONENT+ 2*`MANTISSA + 4:`EXPONENT+ 2*`MANTISSA + 5] CExp_0
[`EXPONENT+ 2*`MANTISSA + 4 : 2*`MANTISSA + 5] Shift_0
[2*`MANTISSA + 4:`MANTISSA + 5] Mmax_0
[`MANTISSA + 4 : `MANTISSA] InputExc_0
[`MANTISSA-1:0] MminS_1
*/
			//pipe_2 <= {pipe_1[2*`EXPONENT + 2*`DWIDTH + 5], pipe_1[2*`EXPONENT +6:2*`EXPONENT +5], MaxAB_1, CExp_1[`EXPONENT-1:0], Shift_1[`EXPONENT-1:0], Mmax_1[`MANTISSA-1:0], pipe_1[4:0], MminS_1[`MANTISSA-1:0]} ;	
/* PIPE_3
[2*`EXPONENT+ 2*`MANTISSA + 9] operation
[2*`EXPONENT+ 2*`MANTISSA + 8] Sa_0
[2*`EXPONENT+ 2*`MANTISSA + 7] Sb_0
[2*`EXPONENT+ 2*`MANTISSA + 6] MaxAB_0
[2*`EXPONENT+ 2*`MANTISSA + 5:`EXPONENT+ 2*`MANTISSA + 6] CExp_0
[`EXPONENT+ 2*`MANTISSA + 5 : 2*`MANTISSA + 6] Shift_0
[2*`MANTISSA + 5:`MANTISSA + 6] Mmax_0
[`MANTISSA + 5 : `MANTISSA + 1] InputExc_0
[`MANTISSA:0] MminS_2
*/
			pipe_3 <= {pipe_2[2*`EXPONENT+ 2*`MANTISSA + 8:`MANTISSA], MminS_2[`MANTISSA:0]} ;	
/* PIPE_4
[2*`EXPONENT+ 2*`MANTISSA + 9] operation
[2*`EXPONENT+ 2*`MANTISSA + 8] Sa_0
[2*`EXPONENT+ 2*`MANTISSA + 7] Sb_0
[2*`EXPONENT+ 2*`MANTISSA + 6] MaxAB_0
[2*`EXPONENT+ 2*`MANTISSA + 5:`EXPONENT+ 2*`MANTISSA + 6] CExp_0
[`EXPONENT+ 2*`MANTISSA + 5 : 2*`MANTISSA + 6] Shift_0
[2*`MANTISSA + 5:`MANTISSA + 6] Mmax_0
[`MANTISSA + 5 : `MANTISSA + 1] InputExc_0
[`MANTISSA:0] MminS_3
*/				
			//pipe_4 <= {pipe_3[2*`EXPONENT+ 2*`MANTISSA + 9:`MANTISSA+1], Mmin_3[`MANTISSA:0]} ;	
/* PIPE_5 :
[`DWIDTH+ `EXPONENT + 11] operation
[`DWIDTH+ `EXPONENT + 10] PSgn_4
[`DWIDTH+ `EXPONENT + 9] Opr_4
[`DWIDTH+ `EXPONENT + 8] Sa_0
[`DWIDTH+ `EXPONENT + 7] Sb_0
[`DWIDTH+ `EXPONENT + 6] MaxAB_0
[`DWIDTH+ `EXPONENT + 5 :`DWIDTH+6] CExp_0
[`DWIDTH+5:`DWIDTH+1] InputExc_0
[`DWIDTH:0] Sum_4
*/					
			pipe_5 <= {pipe_4[2*`EXPONENT+ 2*`MANTISSA + 9], PSgn_4, Opr_4, pipe_4[2*`EXPONENT+ 2*`MANTISSA + 8:`EXPONENT+ 2*`MANTISSA + 6], pipe_4[`MANTISSA+5:`MANTISSA+1], Sum_4[`DWIDTH:0]} ;
/* PIPE_6 :
[`DWIDTH+ `EXPONENT + 16] operation
[`DWIDTH+ `EXPONENT + 15:`DWIDTH+ `EXPONENT + 11] Shift_5
[`DWIDTH+ `EXPONENT + 10] PSgn_4
[`DWIDTH+ `EXPONENT + 9] Opr_4
[`DWIDTH+ `EXPONENT + 8] Sa_0
[`DWIDTH+ `EXPONENT + 7] Sb_0
[`DWIDTH+ `EXPONENT + 6] MaxAB_0
[`DWIDTH+ `EXPONENT + 5 :`DWIDTH+6] CExp_0
[`DWIDTH+5:`DWIDTH+1] InputExc_0
[`DWIDTH:0] Sum_4
*/				
			//pipe_6 <= {pipe_5[`DWIDTH+`EXPONENT+11], Shift_5[4:0], pipe_5[`DWIDTH+`EXPONENT+10:`DWIDTH+1], SumS_5[`DWIDTH:0]} ;	
/* PIPE_7 :
[`DWIDTH+ `EXPONENT + 16] operation
[`DWIDTH+ `EXPONENT + 15:`DWIDTH+ `EXPONENT + 11] Shift_5
[`DWIDTH+ `EXPONENT + 10] PSgn_4
[`DWIDTH+ `EXPONENT + 9] Opr_4
[`DWIDTH+ `EXPONENT + 8] Sa_0
[`DWIDTH+ `EXPONENT + 7] Sb_0
[`DWIDTH+ `EXPONENT + 6] MaxAB_0
[`DWIDTH+ `EXPONENT + 5 :`DWIDTH+6] CExp_0
[`DWIDTH+5:`DWIDTH+1] InputExc_0
[`DWIDTH:0] Sum_4
*/						
			//pipe_7 <= {pipe_6[`DWIDTH+`EXPONENT+16:`DWIDTH+1], SumS_7[`DWIDTH:0]} ;	
/* PIPE_8:
[2*`EXPONENT + `MANTISSA + 15] FG_8 
[2*`EXPONENT + `MANTISSA + 14] operation
[2*`EXPONENT + `MANTISSA + 13] PSgn_4
[2*`EXPONENT + `MANTISSA + 12] Sa_0
[2*`EXPONENT + `MANTISSA + 11] Sb_0
[2*`EXPONENT + `MANTISSA + 10] MaxAB_0
[2*`EXPONENT + `MANTISSA + 9:`EXPONENT + `MANTISSA + 10] CExp_0
[`EXPONENT + `MANTISSA + 9:`EXPONENT + `MANTISSA + 5] InputExc_8
[`EXPONENT + `MANTISSA + 4 :`EXPONENT + 5] NormM_8 
[`EXPONENT + 4 :4] NormE_8
[3] ZeroSum_8
[2] NegE_8
[1] R_8
[0] S_8
*/				
			pipe_8 <= {FG_8, pipe_7[`DWIDTH+`EXPONENT+16], pipe_7[`DWIDTH+`EXPONENT+10], pipe_7[`DWIDTH+`EXPONENT+8:`DWIDTH+1], NormM_8[`MANTISSA-1:0], NormE_8[`EXPONENT:0], ZeroSum_8, NegE_8, R_8, S_8} ;	
/* pipe_9:
[`DWIDTH + 8 :9] P_int
[8] NegE_8
[7] R_8
[6] S_8
[5:1] InputExc_8
[0] EOF
*/				
			//pipe_9 <= {P_int[`DWIDTH-1:0], pipe_8[2], pipe_8[1], pipe_8[0], pipe_8[`EXPONENT+`MANTISSA+9:`EXPONENT+`MANTISSA+5], EOF} ;	
		end
	end		
	
endmodule


//
// Description:	 	The pre-alignment module is responsible for taking the inputs
//							apart and checking the parts for exceptions.
//							The exponent difference is also calculated in this module.
//


module FPAddSub_PrealignModule(
		A,
		B,
		operation,
		Sa,
		Sb,
		ShiftDet,
		InputExc,
		Aout,
		Bout,
		Opout
	);
	
	// Input ports
	input [`DWIDTH-1:0] A ;										// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	// Output ports
	output Sa ;												// A's sign
	output Sb ;												// B's sign
	output [2*`EXPONENT-1:0] ShiftDet ;
	output [4:0] InputExc ;								// Input numbers are exceptions
	output [`DWIDTH-2:0] Aout ;
	output [`DWIDTH-2:0] Bout ;
	output Opout ;
	
	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [`EXPONENT-1:0] DAB ;										// ExpA - ExpB					
	wire [`EXPONENT-1:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & |(A[`MANTISSA-1:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & |(B[`MANTISSA-1:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & ~|(A[`MANTISSA-1:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & ~|(B[`MANTISSA-1:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
	assign DAB = (A[`DWIDTH-2:`MANTISSA] + ~(B[`DWIDTH-2:`MANTISSA]) + 1) ;
	assign DBA = (B[`DWIDTH-2:`MANTISSA] + ~(A[`DWIDTH-2:`MANTISSA]) + 1) ;
	
	assign Sa = A[`DWIDTH-1] ;									// A's sign bit
	assign Sb = B[`DWIDTH-1] ;									// B's sign	bit
	assign ShiftDet = {DBA[`EXPONENT-1:0], DAB[`EXPONENT-1:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[`DWIDTH-2:0] ;
	assign Bout = B[`DWIDTH-2:0] ;
	
endmodule


//
// Description:	 	The alignment module determines the larger input operand and
//							sets the mantissas, shift and common exponent accordingly.
//


module FPAddSub_AlignModule (
		A,
		B,
		ShiftDet,
		CExp,
		MaxAB,
		Shift,
		Mmin,
		Mmax
	);
	
	// Input ports
	input [`DWIDTH-2:0] A ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-2:0] B ;								// Input B, a 32-bit floating point number
	input [2*`EXPONENT-1:0] ShiftDet ;
	
	// Output ports
	output [`EXPONENT-1:0] CExp ;							// Common Exponent
	output MaxAB ;									// Incidates larger of A and B (0/A, 1/B)
	output [`EXPONENT-1:0] Shift ;							// Number of steps to smaller mantissa shift right
	output [`MANTISSA-1:0] Mmin ;							// Smaller mantissa 
	output [`MANTISSA-1:0] Mmax ;							// Larger mantissa
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (A[`DWIDTH-2:0] < B[`DWIDTH-2:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[2*`EXPONENT-1:`EXPONENT] : ShiftDet[`EXPONENT-1:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin = MaxAB ? A[`MANTISSA-1:0] : B[`MANTISSA-1:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? B[`MANTISSA-1:0]: A[`MANTISSA-1:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? B[`MANTISSA+`EXPONENT-1:`MANTISSA] : A[`MANTISSA+`EXPONENT-1:`MANTISSA]) ;		
	
endmodule


// Description:	 Alignment shift stage 1, performs 16|12|8|4 shift
//


// ONLY THIS MODULE IS HARDCODED for half precision fp16 and bfloat16
module FPAddSub_AlignShift1(
		//bf16,
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	//input bf16;
	input [`MANTISSA-1:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [`EXPONENT-3:0] Shift ;						// Shift amount. Last 2 bits of shifting are done in next stage. Hence, we have [`EXPONENT - 2] bits
	
	// Output ports
	output [`MANTISSA:0] Mmin ;						// The smaller mantissa
	

	wire bf16;
	assign bf16 = 1'b1; //hardcoding to 1, to avoid ODIN issue. a `ifdef here wasn't working. apparently, nested `ifdefs don't work

	// Internal signals
	reg	  [`MANTISSA:0]		Lvl1;
	reg	  [`MANTISSA:0]		Lvl2;
	wire    [2*`MANTISSA+1:0]    Stage1;	
	integer           i;                // Loop variable

	wire [`MANTISSA:0] temp_0; 

assign temp_0 = 0;

	always @(*) begin
		if (bf16 == 1'b1) begin						
//hardcoding for bfloat16
	//For bfloat16, we can shift the mantissa by a max of 7 bits since mantissa has a width of 7. 
	//Hence if either, bit[3]/bit[4]/bit[5]/bit[6]/bit[7] is 1, we can make it 0. This corresponds to bits [5:1] in our updated shift which doesn't contain last 2 bits.
		//Lvl1 <= (Shift[1]|Shift[2]|Shift[3]|Shift[4]|Shift[5]) ? {temp_0} : {1'b1, MminP};  // MANTISSA + 1 width	
		Lvl1 <= (|Shift[`EXPONENT-3:1]) ? {temp_0} : {1'b1, MminP};  // MANTISSA + 1 width	
		end
		else begin
		//for half precision fp16, 10 bits can be shifted. Hence, only shifts till 10 (01010)can be made. 
		Lvl1 <= Shift[2] ? {temp_0} : {1'b1, MminP};
		end
	end
	
	assign Stage1 = { temp_0, Lvl1}; //2*MANTISSA + 2 width

	always @(*) begin    					// Rotate {0 | 4 } bits
	if(bf16 == 1'b1) begin
	  case (Shift[0])
			// Rotate by 0	
			1'b0:  Lvl2 <= Stage1[`MANTISSA:0];       			
			// Rotate by 4	
			1'b1:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[`MANTISSA:`MANTISSA-3] <= 0; end
	  endcase
	end
	else begin
	  case (Shift[1:0])					// Rotate {0 | 4 | 8} bits
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[`MANTISSA:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[`MANTISSA:`MANTISSA-3] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[`MANTISSA:`MANTISSA-7] <= 0; end
			// Rotate by 12	
			2'b11: Lvl2[`MANTISSA: 0] <= 0; 
			//2'b11:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[`MANTISSA:`MANTISSA-12] <= 0; end
	  endcase
	end
	end

	// Assign output to next shift stage
	assign Mmin = Lvl2;
	
endmodule


// Description:	 Alignment shift stage 2, performs 3|2|1 shift
//


module FPAddSub_AlignShift2(
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	input [`MANTISSA:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [1:0] Shift ;						// Shift amount. Last 2 bits
	
	// Output ports
	output [`MANTISSA:0] Mmin ;						// The smaller mantissa
	
	// Internal Signal
	reg	  [`MANTISSA:0]		Lvl3;
	wire    [2*`MANTISSA+1:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {11'b0, MminP};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[`MANTISSA:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[`MANTISSA] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[`MANTISSA:`MANTISSA-1] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[`MANTISSA:`MANTISSA-2] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin = Lvl3;						// Take out smaller mantissa				

endmodule


//
// Description:	 Module that executes the addition or subtraction on mantissas.
//


module FPAddSub_ExecutionModule(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		Sum,
		PSgn,
		Opr
    );

	// Input ports
	input [`MANTISSA-1:0] Mmax ;					// The larger mantissa
	input [`MANTISSA:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	output [`DWIDTH:0] Sum ;					// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	wire [`EXPONENT-1:0]temp_1;

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation
	assign temp_1 = 0;
	// Perform effective operation
//SAMIDH_UNSURE 5--> 8

	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, temp_1} - {Mmin, temp_1}) : ({1'b1, Mmax, temp_1} + {Mmin, temp_1}) ;
	
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

endmodule


//
// Description:	 Determine the normalization shift amount and perform 16-shift
//


module FPAddSub_NormalizeModule(
		Sum,
		Mmin,
		Shift
    );

	// Input ports
	input [`DWIDTH:0] Sum ;					// Mantissa sum including hidden 1 and GRS
	
	// Output ports
	output [`DWIDTH:0] Mmin ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount
	//Changes in this doesn't matter since even Bfloat16 can't go beyond 7 shift to the mantissa (only 3 bits valid here)  
	// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[16] ? 5'b00000 :	 
		Sum[15] ? 5'b00001 : 
		Sum[14] ? 5'b00010 : 
		Sum[13] ? 5'b00011 : 
		Sum[12] ? 5'b00100 : 
		Sum[11] ? 5'b00101 : 
		Sum[10] ? 5'b00110 : 
		Sum[9] ? 5'b00111 :
		Sum[8] ? 5'b01000 :
		Sum[7] ? 5'b01001 :
		Sum[6] ? 5'b01010 :
		Sum[5] ? 5'b01011 :
		Sum[4] ? 5'b01100 : 5'b01101
	//	Sum[19] ? 5'b01101 :
	//	Sum[18] ? 5'b01110 :
	//	Sum[17] ? 5'b01111 :
	//	Sum[16] ? 5'b10000 :
	//	Sum[15] ? 5'b10001 :
	//	Sum[14] ? 5'b10010 :
	//	Sum[13] ? 5'b10011 :
	//	Sum[12] ? 5'b10100 :
	//	Sum[11] ? 5'b10101 :
	//	Sum[10] ? 5'b10110 :
	//	Sum[9] ? 5'b10111 :
	//	Sum[8] ? 5'b11000 :
	//	Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [`DWIDTH:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[8:0], 8'b00000000} : Sum; 
	end
	
	// Assign outputs
	assign Mmin = Lvl1;						// Take out smaller mantissa

endmodule


// Description:	 Normalization shift stage 1, performs 12|8|4|3|2|1|0 shift
//
//Hardcoding loop start and end values of i. To avoid ODIN limitations. i=`DWIDTH*2+1 wasn't working.

module FPAddSub_NormalizeShift1(
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	input [`DWIDTH:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [3:0] Shift ;						// Shift amount
	
	// Output ports
	output [`DWIDTH:0] Mmin ;						// The smaller mantissa
	
	reg	  [`DWIDTH:0]		Lvl2;
	wire    [2*`DWIDTH+1:0]    Stage1;	
	reg	  [`DWIDTH:0]		Lvl3;
	wire    [2*`DWIDTH+1:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {MminP, MminP};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[`DWIDTH:0];       		
			// Rotate by 4
			2'b01: begin for (i=33; i>=17; i=i-1) begin Lvl2[i-`DWIDTH -1] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=33; i>=17; i=i-1) begin Lvl2[i-`DWIDTH -1] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=33; i>=17; i=i-1) begin Lvl2[i-`DWIDTH -1] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[`DWIDTH:0];
			// Rotate by 1
			2'b01: begin for (i=33; i>=17; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=33; i>=17; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=33; i>=17; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign Mmin = Lvl3;						// Take out smaller mantissa			
	
endmodule


// Description:	 Normalization shift stage 2, calculates post-normalization
//						 mantissa and exponent, as well as the bits used in rounding		
//


module FPAddSub_NormalizeShift2(
		PSSum,
		CExp,
		Shift,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [`DWIDTH:0] PSSum ;					// The Pre-Shift-Sum
	input [`EXPONENT-1:0] CExp ;
	input [4:0] Shift ;					// Amount to be shifted

	// Output ports
	output [`MANTISSA-1:0] NormM ;				// Normalized mantissa
	output [`EXPONENT:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;

	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [`EXPONENT:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [`EXPONENT:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = PSSum[`DWIDTH] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|PSSum ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[`EXPONENT] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = PSSum[`DWIDTH-1:`EXPONENT+1] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = PSSum[`EXPONENT] ; 
	assign R = PSSum[`EXPONENT-1] ;
	assign S = |PSSum[`EXPONENT-2:0] ;
	
endmodule


// Description:	 Performs 'Round to nearest, tie to even'-rounding on the
//						 normalized mantissa according to the G, R, S bits. Calculates
//						 final result and checks for exponent overflow.
//


module FPAddSub_RoundModule(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		Z,
		EOF
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [`EXPONENT:0] NormE ;				// Normalized exponent
	input [`MANTISSA-1:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	
	// Output ports
	output [`DWIDTH-1:0] Z ;					// Final result
	output EOF ;
	
	// Internal signals
	wire [`MANTISSA:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [`MANTISSA-1:0] RoundM ;				// The final rounded sum
	wire [`EXPONENT:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
        wire FSgn;
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	
	wire [`EXPONENT:0]temp_2;
	assign temp_2 = 0;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[`MANTISSA-1:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[`MANTISSA] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? temp_2 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[`EXPONENT-1:0], RoundM[`MANTISSA-1:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[`EXPONENT];
	
endmodule


//
// Description:	 Check the final result for exception conditions and set
//						 flags accordingly.
//


module FPAddSub_ExceptionModule(
		Z,
		NegE,
		R,
		S,
		InputExc,
		EOF,
		P,
		Flags
    );
	 
	// Input ports
	input [`DWIDTH-1:0] Z	;					// Final product
	input NegE ;						// Negative exponent?
	input R ;							// Round bit
	input S ;							// Sticky bit
	input [4:0] InputExc ;			// Exceptions in inputs A and B
	input EOF ;
	
	// Output ports
	output [`DWIDTH-1:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[`MANTISSA+`EXPONENT-1:`MANTISSA]) & ~|(Z[`MANTISSA+`EXPONENT-1:`MANTISSA]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule
module adder_tree_3stage_16bit (clk,reset,inp00,inp01,inp10,inp11,inp20,inp21,inp30,inp31,sum_out); 

input clk; 
input reset; 
input [15:0] inp00; 
input [15:0] inp01;
input [15:0] inp10; 
input [15:0] inp11;
input [15:0] inp20; 
input [15:0] inp21;
input [15:0] inp30; 
input [15:0] inp31;
output reg [31:0] sum_out;

reg [16:0] S_0_0; 
reg [16:0] S_0_1;
reg [16:0] S_0_2;
reg [16:0] S_0_3;

always@(posedge clk) begin 

S_0_0 <= inp00 + inp01; 
S_0_1 <= inp10 + inp11;
S_0_2 <= inp20 + inp21;
S_0_3 <= inp30 + inp31;

end 

reg [17:0] S_1_0;
reg [17:0] S_1_1;

always@(posedge clk) begin 

S_1_0 <= S_0_0 + S_0_1; 
S_1_1 <= S_0_2 + S_0_3;

end 

always@(posedge clk) begin 

if (reset == 1'b1) begin 
  sum_out <= 32'd0; 
end
else begin 
  sum_out <= S_1_0 + S_1_1; 
end

end 

endmodule 
