
module top (input clk, input reset,input [543:0] top_inp, output [1845:0] top_outp); 
 


 wire [415:0] inp_dpram1;
wire [319:0] outp_dpram1;

dpram_2048_40bit_module_4 dpram1 (.clk(clk),.reset(reset),.inp(inp_dpram1),.outp(outp_dpram1)); 


 wire [2047:0] inp_dsp_ch1;
wire [255:0] outp_dsp_ch1;

dsp_chain_4_fp16_sop2_mult_module_8 dsp_ch1 (.clk(clk),.reset(reset),.inp(inp_dsp_ch1),.outp(outp_dsp_ch1)); 
wire [319:0] inp_interface_1; 
wire [2047:0] outp_interface_1; 

interface_1 inst_interface_1(.clk(clk),.reset(reset),.inp(inp_interface_1),.outp(outp_interface_1)); 


 wire [511:0] inp_dsp_ch2;
wire [127:0] outp_dsp_ch2;

dsp_chain_2_fp16_sop2_mult_module_4 dsp_ch2 (.clk(clk),.reset(reset),.inp(inp_dsp_ch2),.outp(outp_dsp_ch2)); 
wire [319:0] inp_interface_2; 
wire [511:0] outp_interface_2; 

interface_2 inst_interface_2(.clk(clk),.reset(reset),.inp(inp_interface_2),.outp(outp_interface_2)); 


 wire [1151:0] inp_dsp_ch3;
wire [191:0] outp_dsp_ch3;

dsp_chain_3_fp16_sop2_mult_module_6 dsp_ch3 (.clk(clk),.reset(reset),.inp(inp_dsp_ch3),.outp(outp_dsp_ch3)); 
wire [319:0] inp_interface_3; 
wire [1151:0] outp_interface_3; 

interface_3 inst_interface_3(.clk(clk),.reset(reset),.inp(inp_interface_3),.outp(outp_interface_3)); 


 wire [1043:0] inp_activ1;
wire [1031:0] outp_activ1;

activation_32_8bit_module_4 activ1 (.clk(clk),.reset(reset),.inp(inp_activ1),.outp(outp_activ1)); 
wire [255:0] inp_interface_4; 
wire [1043:0] outp_interface_4; 

interface_4 inst_interface_4(.clk(clk),.reset(reset),.inp(inp_interface_4),.outp(outp_interface_4)); 


 wire [1547:0] inp_activ2;
wire [1541:0] outp_activ2;

activation_32_16bit_module_3 activ2 (.clk(clk),.reset(reset),.inp(inp_activ2),.outp(outp_activ2)); 
wire [255:0] inp_interface_5; 
wire [1547:0] outp_interface_5; 

interface_5 inst_interface_5(.clk(clk),.reset(reset),.inp(inp_interface_5),.outp(outp_interface_5)); 


 wire [191:0] inp_activ3;
wire [191:0] outp_activ3;

tanh_16bit_12 activ3 (.clk(clk),.reset(reset),.inp(inp_activ3),.outp(outp_activ3)); 
wire [127:0] inp_interface_6; 
wire [191:0] outp_interface_6; 

interface_6 inst_interface_6(.clk(clk),.reset(reset),.inp(inp_interface_6),.outp(outp_interface_6)); 


 wire [1565:0] inp_activ4;
wire [1547:0] outp_activ4;

activation_32_8bit_module_6 activ4 (.clk(clk),.reset(reset),.inp(inp_activ4),.outp(outp_activ4)); 
wire [127:0] inp_interface_7; 
wire [1565:0] outp_interface_7; 

interface_7 inst_interface_7(.clk(clk),.reset(reset),.inp(inp_interface_7),.outp(outp_interface_7)); 


 wire [383:0] inp_activ5;
wire [383:0] outp_activ5;

sigmoid_16bit_24 activ5 (.clk(clk),.reset(reset),.inp(inp_activ5),.outp(outp_activ5)); 
wire [191:0] inp_interface_8; 
wire [383:0] outp_interface_8; 

interface_8 inst_interface_8(.clk(clk),.reset(reset),.inp(inp_interface_8),.outp(outp_interface_8)); 


 wire [2087:0] inp_activ6;
wire [2063:0] outp_activ6;

activation_32_8bit_module_8 activ6 (.clk(clk),.reset(reset),.inp(inp_activ6),.outp(outp_activ6)); 
wire [191:0] inp_interface_9; 
wire [2087:0] outp_interface_9; 

interface_9 inst_interface_9(.clk(clk),.reset(reset),.inp(inp_interface_9),.outp(outp_interface_9)); 


 wire [1059:0] inp_dpram2;
wire [799:0] outp_dpram2;

dpram_4096_40bit_module_10 dpram2 (.clk(clk),.reset(reset),.inp(inp_dpram2),.outp(outp_dpram2)); 
wire [1031:0] inp_interface_10; 
wire [1059:0] outp_interface_10; 

interface_10 inst_interface_10(.clk(clk),.reset(reset),.inp(inp_interface_10),.outp(outp_interface_10)); 


 wire [1167:0] inp_dpram3;
wire [959:0] outp_dpram3;

dpram_4096_60bit_module_8 dpram3 (.clk(clk),.reset(reset),.inp(inp_dpram3),.outp(outp_dpram3)); 
wire [1541:0] inp_interface_11; 
wire [1167:0] outp_interface_11; 

interface_11 inst_interface_11(.clk(clk),.reset(reset),.inp(inp_interface_11),.outp(outp_interface_11)); 


 wire [2879:0] inp_dpram4;
wire [2399:0] outp_dpram4;

dpram_2048_60bit_module_20 dpram4 (.clk(clk),.reset(reset),.inp(inp_dpram4),.outp(outp_dpram4)); 
wire [191:0] inp_interface_12; 
wire [2879:0] outp_interface_12; 

interface_12 inst_interface_12(.clk(clk),.reset(reset),.inp(inp_interface_12),.outp(outp_interface_12)); 


 wire [2495:0] inp_dpram5;
wire [1919:0] outp_dpram5;

dpram_2048_40bit_module_24 dpram5 (.clk(clk),.reset(reset),.inp(inp_dpram5),.outp(outp_dpram5)); 
wire [1547:0] inp_interface_13; 
wire [2495:0] outp_interface_13; 

interface_13 inst_interface_13(.clk(clk),.reset(reset),.inp(inp_interface_13),.outp(outp_interface_13)); 


 wire [2331:0] inp_dpram6;
wire [1759:0] outp_dpram6;

dpram_4096_40bit_module_22 dpram6 (.clk(clk),.reset(reset),.inp(inp_dpram6),.outp(outp_dpram6)); 
wire [383:0] inp_interface_14; 
wire [2331:0] outp_interface_14; 

interface_14 inst_interface_14(.clk(clk),.reset(reset),.inp(inp_interface_14),.outp(outp_interface_14)); 


 wire [4319:0] inp_dpram7;
wire [3599:0] outp_dpram7;

dpram_2048_60bit_module_30 dpram7 (.clk(clk),.reset(reset),.inp(inp_dpram7),.outp(outp_dpram7)); 
wire [2063:0] inp_interface_15; 
wire [4319:0] outp_interface_15; 

interface_15 inst_interface_15(.clk(clk),.reset(reset),.inp(inp_interface_15),.outp(outp_interface_15)); 


 wire [127:0] inp_dsp_ch5;
wire [31:0] outp_dsp_ch5;

dsp_chain_2_fp16_sop2_mult_module_1 dsp_ch5 (.clk(clk),.reset(reset),.inp(inp_dsp_ch5),.outp(outp_dsp_ch5)); 


 wire [1695:0] inp_dpram8;
wire [1279:0] outp_dpram8;

dpram_4096_40bit_module_16 dpram8 (.clk(clk),.reset(reset),.inp(inp_dpram8),.outp(outp_dpram8)); 
wire [31:0] inp_interface_17; 
wire [1695:0] outp_interface_17; 

interface_17 inst_interface_17(.clk(clk),.reset(reset),.inp(inp_interface_17),.outp(outp_interface_17)); 


 wire [5119:0] inp_dsp_ch4;
wire [639:0] outp_dsp_ch4;

dsp_chain_4_fp16_sop2_mult_module_20 dsp_ch4 (.clk(clk),.reset(reset),.inp(inp_dsp_ch4),.outp(outp_dsp_ch4)); 
wire [1759:0] inp_interface_18; 
wire [5119:0] outp_interface_18; 

interface_18 inst_interface_18(.clk(clk),.reset(reset),.inp(inp_interface_18),.outp(outp_interface_18)); 


 wire [479:0] inp_activ7;
wire [479:0] outp_activ7;

sigmoid_16bit_30 activ7 (.clk(clk),.reset(reset),.inp(inp_activ7),.outp(outp_activ7)); 
wire [1919:0] inp_interface_19; 
wire [479:0] outp_interface_19; 

interface_19 inst_interface_19(.clk(clk),.reset(reset),.inp(inp_interface_19),.outp(outp_interface_19)); 


 wire [4991:0] inp_dsp_ch6;
wire [831:0] outp_dsp_ch6;

dsp_chain_3_fp16_sop2_mult_module_26 dsp_ch6 (.clk(clk),.reset(reset),.inp(inp_dsp_ch6),.outp(outp_dsp_ch6)); 
wire [6079:0] inp_interface_20; 
wire [4991:0] outp_interface_20; 

interface_20 inst_interface_20(.clk(clk),.reset(reset),.inp(inp_interface_20),.outp(outp_interface_20)); 


 wire [2063:0] inp_activ8;
wire [2055:0] outp_activ8;

activation_32_16bit_module_4 activ8 (.clk(clk),.reset(reset),.inp(inp_activ8),.outp(outp_activ8)); 
wire [831:0] inp_interface_21; 
wire [2063:0] outp_interface_21; 

interface_21 inst_interface_21(.clk(clk),.reset(reset),.inp(inp_interface_21),.outp(outp_interface_21)); 


 wire [311:0] inp_dpram9;
wire [239:0] outp_dpram9;

dpram_2048_40bit_module_3 dpram9 (.clk(clk),.reset(reset),.inp(inp_dpram9),.outp(outp_dpram9)); 
wire [2055:0] inp_interface_22; 
wire [311:0] outp_interface_22; 

interface_22 inst_interface_22(.clk(clk),.reset(reset),.inp(inp_interface_22),.outp(outp_interface_22)); 


 wire [9599:0] inp_dsp_ch7;
wire [1599:0] outp_dsp_ch7;

dsp_chain_3_fp16_sop2_mult_module_50 dsp_ch7 (.clk(clk),.reset(reset),.inp(inp_dsp_ch7),.outp(outp_dsp_ch7)); 
wire [9679:0] inp_interface_23; 
wire [9599:0] outp_interface_23; 

interface_23 inst_interface_23(.clk(clk),.reset(reset),.inp(inp_interface_23),.outp(outp_interface_23)); 


 wire [5119:0] inp_dsp_ch8;
wire [639:0] outp_dsp_ch8;

dsp_chain_4_fp16_sop2_mult_module_20 dsp_ch8 (.clk(clk),.reset(reset),.inp(inp_dsp_ch8),.outp(outp_dsp_ch8)); 
wire [4319:0] inp_interface_24; 
wire [5119:0] outp_interface_24; 

interface_24 inst_interface_24(.clk(clk),.reset(reset),.inp(inp_interface_24),.outp(outp_interface_24)); 


 wire [527:0] inp_adder_tree1;
wire [63:0] outp_adder_tree1;

adder_tree_3_fp16bit_4 adder_tree1 (.clk(clk),.reset(reset),.inp(inp_adder_tree1),.outp(outp_adder_tree1)); 
wire [2239:0] inp_interface_25; 
wire [527:0] outp_interface_25; 

interface_25 inst_interface_25(.clk(clk),.reset(reset),.inp(inp_interface_25),.outp(outp_interface_25)); 


 wire [4319:0] inp_dpram10;
wire [3599:0] outp_dpram10;

dpram_2048_60bit_module_30 dpram10 (.clk(clk),.reset(reset),.inp(inp_dpram10),.outp(outp_dpram10)); 
wire [5359:0] inp_interface_26; 
wire [4319:0] outp_interface_26; 

interface_26 inst_interface_26(.clk(clk),.reset(reset),.inp(inp_interface_26),.outp(outp_interface_26)); 


 wire [1547:0] inp_activ9;
wire [1541:0] outp_activ9;

activation_32_16bit_module_3 activ9 (.clk(clk),.reset(reset),.inp(inp_activ9),.outp(outp_activ9)); 
wire [3599:0] inp_interface_27; 
wire [1547:0] outp_interface_27; 

interface_27 inst_interface_27(.clk(clk),.reset(reset),.inp(inp_interface_27),.outp(outp_interface_27)); 

assign inp_dpram1 = top_inp[415:0]; 

assign inp_dsp_ch1 = outp_interface_1; 
assign inp_interface_1 = {outp_dpram1}; 
 

assign inp_dsp_ch2 = outp_interface_2; 
assign inp_interface_2 = {outp_dpram1}; 
 

assign inp_dsp_ch3 = outp_interface_3; 
assign inp_interface_3 = {outp_dpram1}; 
 

assign inp_activ1 = outp_interface_4; 
assign inp_interface_4 = {outp_dsp_ch1}; 
 

assign inp_activ2 = outp_interface_5; 
assign inp_interface_5 = {outp_dsp_ch1}; 
 

assign inp_activ3 = outp_interface_6; 
assign inp_interface_6 = {outp_dsp_ch2}; 
 

assign inp_activ4 = outp_interface_7; 
assign inp_interface_7 = {outp_dsp_ch2}; 
 

assign inp_activ5 = outp_interface_8; 
assign inp_interface_8 = {outp_dsp_ch3}; 
 

assign inp_activ6 = outp_interface_9; 
assign inp_interface_9 = {outp_dsp_ch3}; 
 

assign inp_dpram2 = outp_interface_10; 
assign inp_interface_10 = {outp_activ1}; 
 

assign inp_dpram3 = outp_interface_11; 
assign inp_interface_11 = {outp_activ2}; 
 

assign inp_dpram4 = outp_interface_12; 
assign inp_interface_12 = {outp_activ3}; 
 

assign inp_dpram5 = outp_interface_13; 
assign inp_interface_13 = {outp_activ4}; 
 

assign inp_dpram6 = outp_interface_14; 
assign inp_interface_14 = {outp_activ5}; 
 

assign inp_dpram7 = outp_interface_15; 
assign inp_interface_15 = {outp_activ6}; 
 

assign inp_dsp_ch5 = top_inp[543:416]; 

assign inp_dpram8 = outp_interface_17; 
assign inp_interface_17 = {outp_dsp_ch5}; 
 

assign inp_dsp_ch4 = outp_interface_18; 
assign inp_interface_18 = {outp_dpram2,outp_dpram3}; 
 

assign inp_activ7 = outp_interface_19; 
assign inp_interface_19 = {outp_dsp_ch4,outp_dpram8}; 
 

assign inp_dsp_ch6 = outp_interface_20; 
assign inp_interface_20 = {outp_dpram8,outp_activ7,outp_dpram4,outp_dpram5}; 
 

assign inp_activ8 = outp_interface_21; 
assign inp_interface_21 = {outp_dsp_ch6}; 
 

assign inp_dpram9 = outp_interface_22; 
assign top_outp[239:0] = outp_dpram9; 
assign inp_interface_22 = {outp_activ8}; 
 

assign inp_dsp_ch7 = outp_interface_23; 
assign inp_interface_23 = {outp_dpram6,outp_dpram7,outp_dpram4,outp_dpram5}; 
 

assign inp_dsp_ch8 = outp_interface_24; 
assign inp_interface_24 = {outp_dpram5,outp_dpram4}; 
 

assign inp_adder_tree1 = outp_interface_25; 
assign top_outp[303:240] = outp_adder_tree1; 
assign inp_interface_25 = {outp_dsp_ch7,outp_dsp_ch8}; 
 

assign inp_dpram10 = outp_interface_26; 
assign inp_interface_26 = {outp_dpram6,outp_dpram7}; 
 

assign inp_activ9 = outp_interface_27; 
assign top_outp[1845:304] = outp_activ9; 
assign inp_interface_27 = {outp_dpram10}; 
 

 endmodule 


module interface_1(input reg [319:0] inp, output reg [2047:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[319:0] <= inp ; 
outp[639:320] <= inp ; 
outp[959:640] <= inp ; 
outp[1279:960] <= inp ; 
outp[1599:1280] <= inp ; 
outp[1919:1600] <= inp ; 
outp[2047:1920] <= inp[127:0] ; 
end 
endmodule 

module interface_2(input reg [319:0] inp, output reg [511:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[319:0] <= inp ; 
outp[511:320] <= inp[191:0] ; 
end 
endmodule 

module interface_3(input reg [319:0] inp, output reg [1151:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[319:0] <= inp ; 
outp[639:320] <= inp ; 
outp[959:640] <= inp ; 
outp[1151:960] <= inp[191:0] ; 
end 
endmodule 

module interface_4(input reg [255:0] inp, output reg [1043:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[255:0] <= inp ; 
outp[511:256] <= inp ; 
outp[767:512] <= inp ; 
outp[1023:768] <= inp ; 
outp[1043:1024] <= inp[19:0] ; 
end 
endmodule 

module interface_5(input reg [255:0] inp, output reg [1547:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[255:0] <= inp ; 
outp[511:256] <= inp ; 
outp[767:512] <= inp ; 
outp[1023:768] <= inp ; 
outp[1279:1024] <= inp ; 
outp[1535:1280] <= inp ; 
outp[1547:1536] <= inp[11:0] ; 
end 
endmodule 

module interface_6(input reg [127:0] inp, output reg [191:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[127:0] <= inp ; 
outp[191:128] <= inp[63:0] ; 
end 
endmodule 

module interface_7(input reg [127:0] inp, output reg [1565:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[127:0] <= inp ; 
outp[255:128] <= inp ; 
outp[383:256] <= inp ; 
outp[511:384] <= inp ; 
outp[639:512] <= inp ; 
outp[767:640] <= inp ; 
outp[895:768] <= inp ; 
outp[1023:896] <= inp ; 
outp[1151:1024] <= inp ; 
outp[1279:1152] <= inp ; 
outp[1407:1280] <= inp ; 
outp[1535:1408] <= inp ; 
outp[1565:1536] <= inp[29:0] ; 
end 
endmodule 

module interface_8(input reg [191:0] inp, output reg [383:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[191:0] <= inp ; 
outp[383:192] <= inp ; 
end 
endmodule 

module interface_9(input reg [191:0] inp, output reg [2087:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[191:0] <= inp ; 
outp[383:192] <= inp ; 
outp[575:384] <= inp ; 
outp[767:576] <= inp ; 
outp[959:768] <= inp ; 
outp[1151:960] <= inp ; 
outp[1343:1152] <= inp ; 
outp[1535:1344] <= inp ; 
outp[1727:1536] <= inp ; 
outp[1919:1728] <= inp ; 
outp[2087:1920] <= inp[167:0] ; 
end 
endmodule 

module interface_10(input reg [1031:0] inp, output reg [1059:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[1031:0] <= inp ; 
outp[1059:1032] <= inp[27:0] ; 
end 
endmodule 

module interface_11(input reg [1541:0] inp, output reg [1167:0] outp, input clk, input reset);
reg [1541:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [770:0]intermediate_reg_1; 
 
fsm fsm_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
fsm fsm_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
fsm fsm_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
fsm fsm_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
fsm fsm_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
mux_module mux_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
fsm fsm_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
fsm fsm_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
mux_module mux_module_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
mux_module mux_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
fsm fsm_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
fsm fsm_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
fsm fsm_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
mux_module mux_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
fsm fsm_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
fsm fsm_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
fsm fsm_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
mux_module mux_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
fsm fsm_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
fsm fsm_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
fsm fsm_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
fsm fsm_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
mux_module mux_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
fsm fsm_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
fsm fsm_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
fsm fsm_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
fsm fsm_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
fsm fsm_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
mux_module mux_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
fsm fsm_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
mux_module mux_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
fsm fsm_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
fsm fsm_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
fsm fsm_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
fsm fsm_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
mux_module mux_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
mux_module mux_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
fsm fsm_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
fsm fsm_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
mux_module mux_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
fsm fsm_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
mux_module mux_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
fsm fsm_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
fsm fsm_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
fsm fsm_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
fsm fsm_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
fsm fsm_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
fsm fsm_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
mux_module mux_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
fsm fsm_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
fsm fsm_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
fsm fsm_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
mux_module mux_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
mux_module mux_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
mux_module mux_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
fsm fsm_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
fsm fsm_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
mux_module mux_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
fsm fsm_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
fsm fsm_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
fsm fsm_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
fsm fsm_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
mux_module mux_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
fsm fsm_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
fsm fsm_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
fsm fsm_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
fsm fsm_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
fsm fsm_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
fsm fsm_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
mux_module mux_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
mux_module mux_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
fsm fsm_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
fsm fsm_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
fsm fsm_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
fsm fsm_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
fsm fsm_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
fsm fsm_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
fsm fsm_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
fsm fsm_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
fsm fsm_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
fsm fsm_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
mux_module mux_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
fsm fsm_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
mux_module mux_module_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
mux_module mux_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
fsm fsm_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
fsm fsm_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
fsm fsm_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
mux_module mux_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
fsm fsm_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
mux_module mux_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
fsm fsm_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
fsm fsm_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
fsm fsm_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
fsm fsm_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
fsm fsm_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
fsm fsm_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
mux_module mux_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
fsm fsm_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
fsm fsm_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
mux_module mux_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
fsm fsm_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
mux_module mux_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
fsm fsm_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352])); 
fsm fsm_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
fsm fsm_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
mux_module mux_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
fsm fsm_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
fsm fsm_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
mux_module mux_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
mux_module mux_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
fsm fsm_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
mux_module mux_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
mux_module mux_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
fsm fsm_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
mux_module mux_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
mux_module mux_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
fsm fsm_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
fsm fsm_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
mux_module mux_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
fsm fsm_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
fsm fsm_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
mux_module mux_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
fsm fsm_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
fsm fsm_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
mux_module mux_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
fsm fsm_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
fsm fsm_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
mux_module mux_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
mux_module mux_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
mux_module mux_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
fsm fsm_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
fsm fsm_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
mux_module mux_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
mux_module mux_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
mux_module mux_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
fsm fsm_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
fsm fsm_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
fsm fsm_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
mux_module mux_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
mux_module mux_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
fsm fsm_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
mux_module mux_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
fsm fsm_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
fsm fsm_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
mux_module mux_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
mux_module mux_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
mux_module mux_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
fsm fsm_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
fsm fsm_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
fsm fsm_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
fsm fsm_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
fsm fsm_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
mux_module mux_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
fsm fsm_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
fsm fsm_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
fsm fsm_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
fsm fsm_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
mux_module mux_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
mux_module mux_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
fsm fsm_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
fsm fsm_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
fsm fsm_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
fsm fsm_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
fsm fsm_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
mux_module mux_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
mux_module mux_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
fsm fsm_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
mux_module mux_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
mux_module mux_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
mux_module mux_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
mux_module mux_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
fsm fsm_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
fsm fsm_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
mux_module mux_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
fsm fsm_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
mux_module mux_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
fsm fsm_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
mux_module mux_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
fsm fsm_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
fsm fsm_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
fsm fsm_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
fsm fsm_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
mux_module mux_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
fsm fsm_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
fsm fsm_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
fsm fsm_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
fsm fsm_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
fsm fsm_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
fsm fsm_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
mux_module mux_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
mux_module mux_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
fsm fsm_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
fsm fsm_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
fsm fsm_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
mux_module mux_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
wire [769:0]intermediate_wire_2; 
assign intermediate_wire_2[769] = intermediate_reg_1[770]^intermediate_reg_1[769] ; 
assign intermediate_wire_2[768:0] = intermediate_reg_1[768:0] ; 
always@(posedge clk) begin 
outp [769:0] <= intermediate_wire_2; 
outp[1167:770] <= intermediate_wire_2[397:0] ; 
end 
endmodule 
 

module interface_12(input reg [191:0] inp, output reg [2879:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[191:0] <= inp ; 
outp[383:192] <= inp ; 
outp[575:384] <= inp ; 
outp[767:576] <= inp ; 
outp[959:768] <= inp ; 
outp[1151:960] <= inp ; 
outp[1343:1152] <= inp ; 
outp[1535:1344] <= inp ; 
outp[1727:1536] <= inp ; 
outp[1919:1728] <= inp ; 
outp[2111:1920] <= inp ; 
outp[2303:2112] <= inp ; 
outp[2495:2304] <= inp ; 
outp[2687:2496] <= inp ; 
outp[2879:2688] <= inp ; 
end 
endmodule 

module interface_13(input reg [1547:0] inp, output reg [2495:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[1547:0] <= inp ; 
outp[2495:1548] <= inp[947:0] ; 
end 
endmodule 

module interface_14(input reg [383:0] inp, output reg [2331:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[383:0] <= inp ; 
outp[767:384] <= inp ; 
outp[1151:768] <= inp ; 
outp[1535:1152] <= inp ; 
outp[1919:1536] <= inp ; 
outp[2303:1920] <= inp ; 
outp[2331:2304] <= inp[27:0] ; 
end 
endmodule 

module interface_15(input reg [2063:0] inp, output reg [4319:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[2063:0] <= inp ; 
outp[4127:2064] <= inp ; 
outp[4319:4128] <= inp[191:0] ; 
end 
endmodule 

module interface_17(input reg [31:0] inp, output reg [1695:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[31:0] <= inp ; 
outp[63:32] <= inp ; 
outp[95:64] <= inp ; 
outp[127:96] <= inp ; 
outp[159:128] <= inp ; 
outp[191:160] <= inp ; 
outp[223:192] <= inp ; 
outp[255:224] <= inp ; 
outp[287:256] <= inp ; 
outp[319:288] <= inp ; 
outp[351:320] <= inp ; 
outp[383:352] <= inp ; 
outp[415:384] <= inp ; 
outp[447:416] <= inp ; 
outp[479:448] <= inp ; 
outp[511:480] <= inp ; 
outp[543:512] <= inp ; 
outp[575:544] <= inp ; 
outp[607:576] <= inp ; 
outp[639:608] <= inp ; 
outp[671:640] <= inp ; 
outp[703:672] <= inp ; 
outp[735:704] <= inp ; 
outp[767:736] <= inp ; 
outp[799:768] <= inp ; 
outp[831:800] <= inp ; 
outp[863:832] <= inp ; 
outp[895:864] <= inp ; 
outp[927:896] <= inp ; 
outp[959:928] <= inp ; 
outp[991:960] <= inp ; 
outp[1023:992] <= inp ; 
outp[1055:1024] <= inp ; 
outp[1087:1056] <= inp ; 
outp[1119:1088] <= inp ; 
outp[1151:1120] <= inp ; 
outp[1183:1152] <= inp ; 
outp[1215:1184] <= inp ; 
outp[1247:1216] <= inp ; 
outp[1279:1248] <= inp ; 
outp[1311:1280] <= inp ; 
outp[1343:1312] <= inp ; 
outp[1375:1344] <= inp ; 
outp[1407:1376] <= inp ; 
outp[1439:1408] <= inp ; 
outp[1471:1440] <= inp ; 
outp[1503:1472] <= inp ; 
outp[1535:1504] <= inp ; 
outp[1567:1536] <= inp ; 
outp[1599:1568] <= inp ; 
outp[1631:1600] <= inp ; 
outp[1663:1632] <= inp ; 
outp[1695:1664] <= inp ; 
end 
endmodule 

module interface_18(input reg [1759:0] inp, output reg [5119:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[1759:0] <= inp ; 
outp[3519:1760] <= inp ; 
outp[5119:3520] <= inp[1599:0] ; 
end 
endmodule 

module interface_19(input reg [1919:0] inp, output reg [479:0] outp, input clk, input reset);
reg [1919:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [959:0]intermediate_reg_1; 
 
fsm fsm_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959])); 
fsm fsm_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
fsm fsm_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
fsm fsm_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
mux_module mux_module_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
mux_module mux_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
fsm fsm_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
fsm fsm_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
fsm fsm_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
fsm fsm_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
fsm fsm_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
fsm fsm_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
fsm fsm_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
mux_module mux_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
fsm fsm_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
mux_module mux_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
fsm fsm_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
fsm fsm_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
mux_module mux_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
fsm fsm_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
mux_module mux_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
mux_module mux_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
mux_module mux_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
fsm fsm_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
fsm fsm_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
fsm fsm_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
mux_module mux_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
fsm fsm_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
fsm fsm_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
mux_module mux_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
fsm fsm_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
fsm fsm_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
mux_module mux_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
fsm fsm_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
fsm fsm_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
mux_module mux_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
fsm fsm_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
fsm fsm_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
fsm fsm_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
fsm fsm_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
fsm fsm_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
mux_module mux_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
mux_module mux_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
fsm fsm_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
fsm fsm_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
fsm fsm_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
mux_module mux_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
fsm fsm_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
fsm fsm_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
fsm fsm_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
fsm fsm_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
fsm fsm_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
fsm fsm_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
fsm fsm_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
mux_module mux_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
fsm fsm_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
fsm fsm_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
fsm fsm_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
fsm fsm_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
fsm fsm_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
fsm fsm_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
fsm fsm_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
mux_module mux_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
fsm fsm_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
mux_module mux_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
fsm fsm_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
fsm fsm_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
fsm fsm_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
mux_module mux_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
fsm fsm_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
fsm fsm_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
fsm fsm_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
fsm fsm_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
mux_module mux_module_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
fsm fsm_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
mux_module mux_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
fsm fsm_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
fsm fsm_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
mux_module mux_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
fsm fsm_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
fsm fsm_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
mux_module mux_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
mux_module mux_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
fsm fsm_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
mux_module mux_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
fsm fsm_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
fsm fsm_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
fsm fsm_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
fsm fsm_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
fsm fsm_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
mux_module mux_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
fsm fsm_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
fsm fsm_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
mux_module mux_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
fsm fsm_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
mux_module mux_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
mux_module mux_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
fsm fsm_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532])); 
mux_module mux_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
fsm fsm_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
fsm fsm_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
fsm fsm_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
fsm fsm_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
mux_module mux_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
mux_module mux_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
fsm fsm_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
fsm fsm_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
fsm fsm_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
mux_module mux_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
fsm fsm_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
fsm fsm_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
mux_module mux_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
fsm fsm_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
fsm fsm_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
fsm fsm_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
fsm fsm_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
mux_module mux_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
fsm fsm_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
fsm fsm_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
fsm fsm_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
fsm fsm_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
fsm fsm_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
fsm fsm_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
fsm fsm_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
fsm fsm_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
fsm fsm_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
fsm fsm_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
fsm fsm_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
fsm fsm_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
fsm fsm_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
fsm fsm_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
fsm fsm_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
fsm fsm_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
mux_module mux_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
fsm fsm_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
mux_module mux_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
fsm fsm_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
mux_module mux_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
fsm fsm_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
fsm fsm_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
fsm fsm_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384])); 
mux_module mux_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
fsm fsm_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
fsm fsm_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
fsm fsm_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
fsm fsm_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
fsm fsm_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
fsm fsm_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
mux_module mux_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
fsm fsm_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
fsm fsm_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
fsm fsm_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
fsm fsm_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359])); 
fsm fsm_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
fsm fsm_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
fsm fsm_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
fsm fsm_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
fsm fsm_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
fsm fsm_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
fsm fsm_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
fsm fsm_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
fsm fsm_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
mux_module mux_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
mux_module mux_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
mux_module mux_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
fsm fsm_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
fsm fsm_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
mux_module mux_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
fsm fsm_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
fsm fsm_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
mux_module mux_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
fsm fsm_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
fsm fsm_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
fsm fsm_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
fsm fsm_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
fsm fsm_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
fsm fsm_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
mux_module mux_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
mux_module mux_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
mux_module mux_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
fsm fsm_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
mux_module mux_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
fsm fsm_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
fsm fsm_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
mux_module mux_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
mux_module mux_module_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
fsm fsm_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
fsm fsm_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
mux_module mux_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
mux_module mux_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
fsm fsm_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
mux_module mux_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
mux_module mux_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
fsm fsm_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
fsm fsm_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
fsm fsm_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
fsm fsm_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
mux_module mux_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
fsm fsm_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
mux_module mux_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
fsm fsm_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
mux_module mux_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
fsm fsm_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
mux_module mux_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
mux_module mux_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
fsm fsm_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
mux_module mux_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
mux_module mux_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170])); 
fsm fsm_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
fsm fsm_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
fsm fsm_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
fsm fsm_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
mux_module mux_module_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
fsm fsm_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
fsm fsm_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
fsm fsm_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
fsm fsm_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
mux_module mux_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
mux_module mux_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
fsm fsm_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
fsm fsm_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
mux_module mux_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
fsm fsm_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
fsm fsm_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
mux_module mux_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
mux_module mux_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
fsm fsm_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
mux_module mux_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
fsm fsm_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
fsm fsm_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
mux_module mux_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
mux_module mux_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
mux_module mux_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
mux_module mux_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
fsm fsm_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
mux_module mux_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
fsm fsm_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100])); 
fsm fsm_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
fsm fsm_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
fsm fsm_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
mux_module mux_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
fsm fsm_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
mux_module mux_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
mux_module mux_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
fsm fsm_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
mux_module mux_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
fsm fsm_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
mux_module mux_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
mux_module mux_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65])); 
mux_module mux_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
fsm fsm_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
fsm fsm_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
mux_module mux_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
mux_module mux_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
fsm fsm_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
fsm fsm_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
fsm fsm_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
fsm fsm_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48])); 
fsm fsm_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
fsm fsm_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
mux_module mux_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
fsm fsm_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
mux_module mux_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
fsm fsm_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
mux_module mux_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
fsm fsm_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
mux_module mux_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
fsm fsm_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
fsm fsm_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
fsm fsm_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
mux_module mux_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
fsm fsm_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
fsm fsm_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
mux_module mux_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
mux_module mux_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
reg [479:0]intermediate_reg_2; 
 
fsm fsm_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
fsm fsm_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478])); 
mux_module mux_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473])); 
fsm fsm_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472])); 
fsm fsm_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471])); 
fsm fsm_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470])); 
mux_module mux_module_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468])); 
mux_module mux_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464])); 
fsm fsm_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463])); 
fsm fsm_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462])); 
mux_module mux_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458])); 
mux_module mux_module_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455])); 
mux_module mux_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453])); 
mux_module mux_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451])); 
fsm fsm_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450])); 
fsm fsm_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449])); 
fsm fsm_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448])); 
mux_module mux_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446])); 
mux_module mux_module_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444])); 
mux_module mux_module_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442])); 
mux_module mux_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437])); 
fsm fsm_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436])); 
fsm fsm_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435])); 
mux_module mux_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433])); 
fsm fsm_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432])); 
fsm fsm_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431])); 
fsm fsm_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430])); 
fsm fsm_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429])); 
fsm fsm_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428])); 
fsm fsm_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427])); 
fsm fsm_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426])); 
mux_module mux_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423])); 
fsm fsm_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422])); 
fsm fsm_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421])); 
fsm fsm_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420])); 
mux_module mux_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416])); 
mux_module mux_module_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413])); 
mux_module mux_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410])); 
fsm fsm_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409])); 
mux_module mux_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406])); 
mux_module mux_module_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402])); 
mux_module mux_module_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399])); 
mux_module mux_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396])); 
mux_module mux_module_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393])); 
fsm fsm_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392])); 
fsm fsm_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391])); 
fsm fsm_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390])); 
mux_module mux_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388])); 
fsm fsm_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387])); 
fsm fsm_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386])); 
mux_module mux_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383])); 
mux_module mux_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
fsm fsm_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
fsm fsm_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379])); 
fsm fsm_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378])); 
fsm fsm_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377])); 
mux_module mux_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375])); 
fsm fsm_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374])); 
fsm fsm_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373])); 
fsm fsm_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372])); 
mux_module mux_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
fsm fsm_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369])); 
fsm fsm_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368])); 
mux_module mux_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366])); 
fsm fsm_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365])); 
fsm fsm_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
mux_module mux_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361])); 
mux_module mux_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
fsm fsm_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
fsm fsm_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357])); 
mux_module mux_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355])); 
fsm fsm_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354])); 
mux_module mux_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351])); 
mux_module mux_module_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349])); 
fsm fsm_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348])); 
mux_module mux_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
mux_module mux_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342])); 
mux_module mux_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339])); 
fsm fsm_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338])); 
mux_module mux_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336])); 
fsm fsm_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
fsm fsm_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334])); 
mux_module mux_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
fsm fsm_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
mux_module mux_module_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326])); 
mux_module mux_module_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323])); 
mux_module mux_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
fsm fsm_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319])); 
fsm fsm_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318])); 
mux_module mux_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316])); 
mux_module mux_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312])); 
mux_module mux_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309])); 
mux_module mux_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305])); 
fsm fsm_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304])); 
fsm fsm_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
mux_module mux_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
mux_module mux_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298])); 
mux_module mux_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
fsm fsm_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
fsm fsm_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294])); 
fsm fsm_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
mux_module mux_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290])); 
mux_module mux_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288])); 
fsm fsm_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287])); 
mux_module mux_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
mux_module mux_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
fsm fsm_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282])); 
fsm fsm_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281])); 
mux_module mux_module_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279])); 
mux_module mux_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277])); 
fsm fsm_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276])); 
mux_module mux_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
fsm fsm_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
fsm fsm_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
mux_module mux_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
fsm fsm_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268])); 
mux_module mux_module_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266])); 
mux_module mux_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264])); 
mux_module mux_module_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
mux_module mux_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257])); 
fsm fsm_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
mux_module mux_module_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
mux_module mux_module_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
fsm fsm_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248])); 
fsm fsm_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247])); 
mux_module mux_module_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
mux_module mux_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243])); 
mux_module mux_module_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
mux_module mux_module_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
fsm fsm_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
fsm fsm_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236])); 
fsm fsm_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235])); 
fsm fsm_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
fsm fsm_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233])); 
fsm fsm_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232])); 
mux_module mux_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226])); 
fsm fsm_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
fsm fsm_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224])); 
fsm fsm_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223])); 
mux_module mux_module_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219])); 
fsm fsm_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
mux_module mux_module_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214])); 
fsm fsm_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
mux_module mux_module_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
mux_module mux_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
mux_module mux_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
mux_module mux_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200])); 
fsm fsm_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
fsm fsm_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198])); 
fsm fsm_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197])); 
mux_module mux_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195])); 
fsm fsm_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194])); 
fsm fsm_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193])); 
fsm fsm_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
mux_module mux_module_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190])); 
mux_module mux_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
fsm fsm_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
mux_module mux_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185])); 
fsm fsm_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
mux_module mux_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182])); 
fsm fsm_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181])); 
fsm fsm_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180])); 
fsm fsm_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179])); 
fsm fsm_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178])); 
mux_module mux_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175])); 
mux_module mux_module_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
fsm fsm_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
fsm fsm_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
mux_module mux_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168])); 
mux_module mux_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166])); 
fsm fsm_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
fsm fsm_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164])); 
fsm fsm_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
mux_module mux_module_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161])); 
fsm fsm_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160])); 
fsm fsm_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
mux_module mux_module_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157])); 
mux_module mux_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153])); 
mux_module mux_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
mux_module mux_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148])); 
mux_module mux_module_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146])); 
fsm fsm_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145])); 
fsm fsm_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144])); 
mux_module mux_module_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140])); 
mux_module mux_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136])); 
mux_module mux_module_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
fsm fsm_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133])); 
mux_module mux_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131])); 
fsm fsm_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130])); 
fsm fsm_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129])); 
mux_module mux_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126])); 
fsm fsm_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
fsm fsm_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124])); 
fsm fsm_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123])); 
fsm fsm_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
mux_module mux_module_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119])); 
fsm fsm_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118])); 
fsm fsm_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117])); 
mux_module mux_module_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
fsm fsm_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111])); 
mux_module mux_module_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
fsm fsm_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
fsm fsm_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107])); 
mux_module mux_module_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102])); 
fsm fsm_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
fsm fsm_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100])); 
mux_module mux_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98])); 
fsm fsm_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
fsm fsm_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96])); 
fsm fsm_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95])); 
mux_module mux_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
fsm fsm_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92])); 
mux_module mux_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
mux_module mux_module_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
fsm fsm_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
mux_module mux_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
fsm fsm_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82])); 
fsm fsm_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81])); 
mux_module mux_module_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
mux_module mux_module_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
fsm fsm_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74])); 
mux_module mux_module_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72])); 
mux_module mux_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
mux_module mux_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68])); 
mux_module mux_module_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
mux_module mux_module_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60])); 
mux_module mux_module_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55])); 
fsm fsm_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54])); 
fsm fsm_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
fsm fsm_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
fsm fsm_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51])); 
mux_module mux_module_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
mux_module mux_module_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47])); 
mux_module mux_module_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44])); 
fsm fsm_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
mux_module mux_module_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
mux_module mux_module_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
fsm fsm_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36])); 
mux_module mux_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33])); 
mux_module mux_module_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
fsm fsm_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
mux_module mux_module_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
mux_module mux_module_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25])); 
fsm fsm_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
mux_module mux_module_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22])); 
mux_module mux_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
fsm fsm_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15])); 
mux_module mux_module_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11])); 
mux_module mux_module_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
fsm fsm_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6])); 
mux_module mux_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
fsm fsm_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3])); 
mux_module mux_module_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
fsm fsm_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0])); 
always@(posedge clk) begin 
outp[479:0] <= intermediate_reg_2 ; 
end 
endmodule 
 

module interface_20(input reg [6079:0] inp, output reg [4991:0] outp, input clk, input reset);
reg [6079:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [3039:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6079]),.i2(intermediate_reg_0[6078]),.o(intermediate_reg_1[3039]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6077]),.i2(intermediate_reg_0[6076]),.o(intermediate_reg_1[3038])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6075]),.i2(intermediate_reg_0[6074]),.o(intermediate_reg_1[3037])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6073]),.i2(intermediate_reg_0[6072]),.o(intermediate_reg_1[3036]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6071]),.i2(intermediate_reg_0[6070]),.o(intermediate_reg_1[3035])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6069]),.i2(intermediate_reg_0[6068]),.o(intermediate_reg_1[3034]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6067]),.i2(intermediate_reg_0[6066]),.o(intermediate_reg_1[3033])); 
mux_module mux_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6065]),.i2(intermediate_reg_0[6064]),.o(intermediate_reg_1[3032]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6063]),.i2(intermediate_reg_0[6062]),.o(intermediate_reg_1[3031]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6061]),.i2(intermediate_reg_0[6060]),.o(intermediate_reg_1[3030]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6059]),.i2(intermediate_reg_0[6058]),.o(intermediate_reg_1[3029]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6057]),.i2(intermediate_reg_0[6056]),.o(intermediate_reg_1[3028])); 
fsm fsm_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6055]),.i2(intermediate_reg_0[6054]),.o(intermediate_reg_1[3027])); 
fsm fsm_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6053]),.i2(intermediate_reg_0[6052]),.o(intermediate_reg_1[3026])); 
fsm fsm_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6051]),.i2(intermediate_reg_0[6050]),.o(intermediate_reg_1[3025])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6049]),.i2(intermediate_reg_0[6048]),.o(intermediate_reg_1[3024]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6047]),.i2(intermediate_reg_0[6046]),.o(intermediate_reg_1[3023])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6045]),.i2(intermediate_reg_0[6044]),.o(intermediate_reg_1[3022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6043]),.i2(intermediate_reg_0[6042]),.o(intermediate_reg_1[3021]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6041]),.i2(intermediate_reg_0[6040]),.o(intermediate_reg_1[3020])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6039]),.i2(intermediate_reg_0[6038]),.o(intermediate_reg_1[3019]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6037]),.i2(intermediate_reg_0[6036]),.o(intermediate_reg_1[3018]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6035]),.i2(intermediate_reg_0[6034]),.o(intermediate_reg_1[3017])); 
fsm fsm_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6033]),.i2(intermediate_reg_0[6032]),.o(intermediate_reg_1[3016])); 
fsm fsm_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6031]),.i2(intermediate_reg_0[6030]),.o(intermediate_reg_1[3015])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6029]),.i2(intermediate_reg_0[6028]),.o(intermediate_reg_1[3014]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6027]),.i2(intermediate_reg_0[6026]),.o(intermediate_reg_1[3013])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6025]),.i2(intermediate_reg_0[6024]),.o(intermediate_reg_1[3012]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6023]),.i2(intermediate_reg_0[6022]),.o(intermediate_reg_1[3011]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6021]),.i2(intermediate_reg_0[6020]),.o(intermediate_reg_1[3010]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6019]),.i2(intermediate_reg_0[6018]),.o(intermediate_reg_1[3009]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6017]),.i2(intermediate_reg_0[6016]),.o(intermediate_reg_1[3008])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6015]),.i2(intermediate_reg_0[6014]),.o(intermediate_reg_1[3007]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6013]),.i2(intermediate_reg_0[6012]),.o(intermediate_reg_1[3006])); 
fsm fsm_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6011]),.i2(intermediate_reg_0[6010]),.o(intermediate_reg_1[3005])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6009]),.i2(intermediate_reg_0[6008]),.o(intermediate_reg_1[3004])); 
fsm fsm_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6007]),.i2(intermediate_reg_0[6006]),.o(intermediate_reg_1[3003])); 
fsm fsm_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6005]),.i2(intermediate_reg_0[6004]),.o(intermediate_reg_1[3002])); 
fsm fsm_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6003]),.i2(intermediate_reg_0[6002]),.o(intermediate_reg_1[3001])); 
fsm fsm_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6001]),.i2(intermediate_reg_0[6000]),.o(intermediate_reg_1[3000])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5999]),.i2(intermediate_reg_0[5998]),.o(intermediate_reg_1[2999])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5997]),.i2(intermediate_reg_0[5996]),.o(intermediate_reg_1[2998])); 
fsm fsm_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5995]),.i2(intermediate_reg_0[5994]),.o(intermediate_reg_1[2997])); 
fsm fsm_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5993]),.i2(intermediate_reg_0[5992]),.o(intermediate_reg_1[2996])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5991]),.i2(intermediate_reg_0[5990]),.o(intermediate_reg_1[2995]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5989]),.i2(intermediate_reg_0[5988]),.o(intermediate_reg_1[2994]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5987]),.i2(intermediate_reg_0[5986]),.o(intermediate_reg_1[2993])); 
fsm fsm_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5985]),.i2(intermediate_reg_0[5984]),.o(intermediate_reg_1[2992])); 
mux_module mux_module_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5983]),.i2(intermediate_reg_0[5982]),.o(intermediate_reg_1[2991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5981]),.i2(intermediate_reg_0[5980]),.o(intermediate_reg_1[2990]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5979]),.i2(intermediate_reg_0[5978]),.o(intermediate_reg_1[2989]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5977]),.i2(intermediate_reg_0[5976]),.o(intermediate_reg_1[2988]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5975]),.i2(intermediate_reg_0[5974]),.o(intermediate_reg_1[2987])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5973]),.i2(intermediate_reg_0[5972]),.o(intermediate_reg_1[2986]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5971]),.i2(intermediate_reg_0[5970]),.o(intermediate_reg_1[2985]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5969]),.i2(intermediate_reg_0[5968]),.o(intermediate_reg_1[2984])); 
fsm fsm_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5967]),.i2(intermediate_reg_0[5966]),.o(intermediate_reg_1[2983])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5965]),.i2(intermediate_reg_0[5964]),.o(intermediate_reg_1[2982]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5963]),.i2(intermediate_reg_0[5962]),.o(intermediate_reg_1[2981]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5961]),.i2(intermediate_reg_0[5960]),.o(intermediate_reg_1[2980])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5959]),.i2(intermediate_reg_0[5958]),.o(intermediate_reg_1[2979])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5957]),.i2(intermediate_reg_0[5956]),.o(intermediate_reg_1[2978]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5955]),.i2(intermediate_reg_0[5954]),.o(intermediate_reg_1[2977])); 
fsm fsm_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5953]),.i2(intermediate_reg_0[5952]),.o(intermediate_reg_1[2976])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5951]),.i2(intermediate_reg_0[5950]),.o(intermediate_reg_1[2975])); 
fsm fsm_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5949]),.i2(intermediate_reg_0[5948]),.o(intermediate_reg_1[2974])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5947]),.i2(intermediate_reg_0[5946]),.o(intermediate_reg_1[2973]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5945]),.i2(intermediate_reg_0[5944]),.o(intermediate_reg_1[2972]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5943]),.i2(intermediate_reg_0[5942]),.o(intermediate_reg_1[2971])); 
mux_module mux_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5941]),.i2(intermediate_reg_0[5940]),.o(intermediate_reg_1[2970]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5939]),.i2(intermediate_reg_0[5938]),.o(intermediate_reg_1[2969]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5937]),.i2(intermediate_reg_0[5936]),.o(intermediate_reg_1[2968]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5935]),.i2(intermediate_reg_0[5934]),.o(intermediate_reg_1[2967])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5933]),.i2(intermediate_reg_0[5932]),.o(intermediate_reg_1[2966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5931]),.i2(intermediate_reg_0[5930]),.o(intermediate_reg_1[2965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5929]),.i2(intermediate_reg_0[5928]),.o(intermediate_reg_1[2964]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5927]),.i2(intermediate_reg_0[5926]),.o(intermediate_reg_1[2963]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5925]),.i2(intermediate_reg_0[5924]),.o(intermediate_reg_1[2962])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5923]),.i2(intermediate_reg_0[5922]),.o(intermediate_reg_1[2961]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5921]),.i2(intermediate_reg_0[5920]),.o(intermediate_reg_1[2960])); 
fsm fsm_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5919]),.i2(intermediate_reg_0[5918]),.o(intermediate_reg_1[2959])); 
mux_module mux_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5917]),.i2(intermediate_reg_0[5916]),.o(intermediate_reg_1[2958]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5915]),.i2(intermediate_reg_0[5914]),.o(intermediate_reg_1[2957]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5913]),.i2(intermediate_reg_0[5912]),.o(intermediate_reg_1[2956]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5911]),.i2(intermediate_reg_0[5910]),.o(intermediate_reg_1[2955]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5909]),.i2(intermediate_reg_0[5908]),.o(intermediate_reg_1[2954]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5907]),.i2(intermediate_reg_0[5906]),.o(intermediate_reg_1[2953])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5905]),.i2(intermediate_reg_0[5904]),.o(intermediate_reg_1[2952])); 
fsm fsm_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5903]),.i2(intermediate_reg_0[5902]),.o(intermediate_reg_1[2951])); 
fsm fsm_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5901]),.i2(intermediate_reg_0[5900]),.o(intermediate_reg_1[2950])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5899]),.i2(intermediate_reg_0[5898]),.o(intermediate_reg_1[2949]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5897]),.i2(intermediate_reg_0[5896]),.o(intermediate_reg_1[2948])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5895]),.i2(intermediate_reg_0[5894]),.o(intermediate_reg_1[2947]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5893]),.i2(intermediate_reg_0[5892]),.o(intermediate_reg_1[2946])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5891]),.i2(intermediate_reg_0[5890]),.o(intermediate_reg_1[2945]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5889]),.i2(intermediate_reg_0[5888]),.o(intermediate_reg_1[2944])); 
fsm fsm_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5887]),.i2(intermediate_reg_0[5886]),.o(intermediate_reg_1[2943])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5885]),.i2(intermediate_reg_0[5884]),.o(intermediate_reg_1[2942]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5883]),.i2(intermediate_reg_0[5882]),.o(intermediate_reg_1[2941])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5881]),.i2(intermediate_reg_0[5880]),.o(intermediate_reg_1[2940]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5879]),.i2(intermediate_reg_0[5878]),.o(intermediate_reg_1[2939])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5877]),.i2(intermediate_reg_0[5876]),.o(intermediate_reg_1[2938])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5875]),.i2(intermediate_reg_0[5874]),.o(intermediate_reg_1[2937]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5873]),.i2(intermediate_reg_0[5872]),.o(intermediate_reg_1[2936]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5871]),.i2(intermediate_reg_0[5870]),.o(intermediate_reg_1[2935])); 
mux_module mux_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5869]),.i2(intermediate_reg_0[5868]),.o(intermediate_reg_1[2934]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5867]),.i2(intermediate_reg_0[5866]),.o(intermediate_reg_1[2933]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5865]),.i2(intermediate_reg_0[5864]),.o(intermediate_reg_1[2932]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5863]),.i2(intermediate_reg_0[5862]),.o(intermediate_reg_1[2931])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5861]),.i2(intermediate_reg_0[5860]),.o(intermediate_reg_1[2930]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5859]),.i2(intermediate_reg_0[5858]),.o(intermediate_reg_1[2929]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5857]),.i2(intermediate_reg_0[5856]),.o(intermediate_reg_1[2928])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5855]),.i2(intermediate_reg_0[5854]),.o(intermediate_reg_1[2927]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5853]),.i2(intermediate_reg_0[5852]),.o(intermediate_reg_1[2926])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5851]),.i2(intermediate_reg_0[5850]),.o(intermediate_reg_1[2925]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5849]),.i2(intermediate_reg_0[5848]),.o(intermediate_reg_1[2924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5847]),.i2(intermediate_reg_0[5846]),.o(intermediate_reg_1[2923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5845]),.i2(intermediate_reg_0[5844]),.o(intermediate_reg_1[2922]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5843]),.i2(intermediate_reg_0[5842]),.o(intermediate_reg_1[2921])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5841]),.i2(intermediate_reg_0[5840]),.o(intermediate_reg_1[2920])); 
fsm fsm_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5839]),.i2(intermediate_reg_0[5838]),.o(intermediate_reg_1[2919])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5837]),.i2(intermediate_reg_0[5836]),.o(intermediate_reg_1[2918]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5835]),.i2(intermediate_reg_0[5834]),.o(intermediate_reg_1[2917])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5833]),.i2(intermediate_reg_0[5832]),.o(intermediate_reg_1[2916]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5831]),.i2(intermediate_reg_0[5830]),.o(intermediate_reg_1[2915])); 
mux_module mux_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5829]),.i2(intermediate_reg_0[5828]),.o(intermediate_reg_1[2914]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5827]),.i2(intermediate_reg_0[5826]),.o(intermediate_reg_1[2913]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5825]),.i2(intermediate_reg_0[5824]),.o(intermediate_reg_1[2912])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5823]),.i2(intermediate_reg_0[5822]),.o(intermediate_reg_1[2911]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5821]),.i2(intermediate_reg_0[5820]),.o(intermediate_reg_1[2910]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5819]),.i2(intermediate_reg_0[5818]),.o(intermediate_reg_1[2909])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5817]),.i2(intermediate_reg_0[5816]),.o(intermediate_reg_1[2908])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5815]),.i2(intermediate_reg_0[5814]),.o(intermediate_reg_1[2907]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5813]),.i2(intermediate_reg_0[5812]),.o(intermediate_reg_1[2906]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5811]),.i2(intermediate_reg_0[5810]),.o(intermediate_reg_1[2905])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5809]),.i2(intermediate_reg_0[5808]),.o(intermediate_reg_1[2904]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5807]),.i2(intermediate_reg_0[5806]),.o(intermediate_reg_1[2903])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5805]),.i2(intermediate_reg_0[5804]),.o(intermediate_reg_1[2902]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5803]),.i2(intermediate_reg_0[5802]),.o(intermediate_reg_1[2901])); 
mux_module mux_module_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5801]),.i2(intermediate_reg_0[5800]),.o(intermediate_reg_1[2900]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5799]),.i2(intermediate_reg_0[5798]),.o(intermediate_reg_1[2899]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5797]),.i2(intermediate_reg_0[5796]),.o(intermediate_reg_1[2898]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5795]),.i2(intermediate_reg_0[5794]),.o(intermediate_reg_1[2897]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5793]),.i2(intermediate_reg_0[5792]),.o(intermediate_reg_1[2896]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5791]),.i2(intermediate_reg_0[5790]),.o(intermediate_reg_1[2895]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5789]),.i2(intermediate_reg_0[5788]),.o(intermediate_reg_1[2894])); 
fsm fsm_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5787]),.i2(intermediate_reg_0[5786]),.o(intermediate_reg_1[2893])); 
fsm fsm_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5785]),.i2(intermediate_reg_0[5784]),.o(intermediate_reg_1[2892])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5783]),.i2(intermediate_reg_0[5782]),.o(intermediate_reg_1[2891]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5781]),.i2(intermediate_reg_0[5780]),.o(intermediate_reg_1[2890])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5779]),.i2(intermediate_reg_0[5778]),.o(intermediate_reg_1[2889]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5777]),.i2(intermediate_reg_0[5776]),.o(intermediate_reg_1[2888]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5775]),.i2(intermediate_reg_0[5774]),.o(intermediate_reg_1[2887]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5773]),.i2(intermediate_reg_0[5772]),.o(intermediate_reg_1[2886])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5771]),.i2(intermediate_reg_0[5770]),.o(intermediate_reg_1[2885]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5769]),.i2(intermediate_reg_0[5768]),.o(intermediate_reg_1[2884]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5767]),.i2(intermediate_reg_0[5766]),.o(intermediate_reg_1[2883]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5765]),.i2(intermediate_reg_0[5764]),.o(intermediate_reg_1[2882])); 
mux_module mux_module_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5763]),.i2(intermediate_reg_0[5762]),.o(intermediate_reg_1[2881]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5761]),.i2(intermediate_reg_0[5760]),.o(intermediate_reg_1[2880])); 
fsm fsm_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5759]),.i2(intermediate_reg_0[5758]),.o(intermediate_reg_1[2879])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5757]),.i2(intermediate_reg_0[5756]),.o(intermediate_reg_1[2878]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5755]),.i2(intermediate_reg_0[5754]),.o(intermediate_reg_1[2877])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5753]),.i2(intermediate_reg_0[5752]),.o(intermediate_reg_1[2876]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5751]),.i2(intermediate_reg_0[5750]),.o(intermediate_reg_1[2875]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5749]),.i2(intermediate_reg_0[5748]),.o(intermediate_reg_1[2874]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5747]),.i2(intermediate_reg_0[5746]),.o(intermediate_reg_1[2873])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5745]),.i2(intermediate_reg_0[5744]),.o(intermediate_reg_1[2872]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5743]),.i2(intermediate_reg_0[5742]),.o(intermediate_reg_1[2871]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5741]),.i2(intermediate_reg_0[5740]),.o(intermediate_reg_1[2870])); 
fsm fsm_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5739]),.i2(intermediate_reg_0[5738]),.o(intermediate_reg_1[2869])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5737]),.i2(intermediate_reg_0[5736]),.o(intermediate_reg_1[2868]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5735]),.i2(intermediate_reg_0[5734]),.o(intermediate_reg_1[2867]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5733]),.i2(intermediate_reg_0[5732]),.o(intermediate_reg_1[2866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5731]),.i2(intermediate_reg_0[5730]),.o(intermediate_reg_1[2865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5729]),.i2(intermediate_reg_0[5728]),.o(intermediate_reg_1[2864]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5727]),.i2(intermediate_reg_0[5726]),.o(intermediate_reg_1[2863]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5725]),.i2(intermediate_reg_0[5724]),.o(intermediate_reg_1[2862])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5723]),.i2(intermediate_reg_0[5722]),.o(intermediate_reg_1[2861])); 
fsm fsm_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5721]),.i2(intermediate_reg_0[5720]),.o(intermediate_reg_1[2860])); 
mux_module mux_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5719]),.i2(intermediate_reg_0[5718]),.o(intermediate_reg_1[2859]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5717]),.i2(intermediate_reg_0[5716]),.o(intermediate_reg_1[2858]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5715]),.i2(intermediate_reg_0[5714]),.o(intermediate_reg_1[2857])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5713]),.i2(intermediate_reg_0[5712]),.o(intermediate_reg_1[2856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5711]),.i2(intermediate_reg_0[5710]),.o(intermediate_reg_1[2855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5709]),.i2(intermediate_reg_0[5708]),.o(intermediate_reg_1[2854]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5707]),.i2(intermediate_reg_0[5706]),.o(intermediate_reg_1[2853])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5705]),.i2(intermediate_reg_0[5704]),.o(intermediate_reg_1[2852]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5703]),.i2(intermediate_reg_0[5702]),.o(intermediate_reg_1[2851])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5701]),.i2(intermediate_reg_0[5700]),.o(intermediate_reg_1[2850]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5699]),.i2(intermediate_reg_0[5698]),.o(intermediate_reg_1[2849])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5697]),.i2(intermediate_reg_0[5696]),.o(intermediate_reg_1[2848]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5695]),.i2(intermediate_reg_0[5694]),.o(intermediate_reg_1[2847])); 
fsm fsm_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5693]),.i2(intermediate_reg_0[5692]),.o(intermediate_reg_1[2846])); 
fsm fsm_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5691]),.i2(intermediate_reg_0[5690]),.o(intermediate_reg_1[2845])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5689]),.i2(intermediate_reg_0[5688]),.o(intermediate_reg_1[2844]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5687]),.i2(intermediate_reg_0[5686]),.o(intermediate_reg_1[2843])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5685]),.i2(intermediate_reg_0[5684]),.o(intermediate_reg_1[2842]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5683]),.i2(intermediate_reg_0[5682]),.o(intermediate_reg_1[2841])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5681]),.i2(intermediate_reg_0[5680]),.o(intermediate_reg_1[2840]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5679]),.i2(intermediate_reg_0[5678]),.o(intermediate_reg_1[2839])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5677]),.i2(intermediate_reg_0[5676]),.o(intermediate_reg_1[2838]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5675]),.i2(intermediate_reg_0[5674]),.o(intermediate_reg_1[2837])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5673]),.i2(intermediate_reg_0[5672]),.o(intermediate_reg_1[2836])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5671]),.i2(intermediate_reg_0[5670]),.o(intermediate_reg_1[2835]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5669]),.i2(intermediate_reg_0[5668]),.o(intermediate_reg_1[2834]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5667]),.i2(intermediate_reg_0[5666]),.o(intermediate_reg_1[2833])); 
mux_module mux_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5665]),.i2(intermediate_reg_0[5664]),.o(intermediate_reg_1[2832]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5663]),.i2(intermediate_reg_0[5662]),.o(intermediate_reg_1[2831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5661]),.i2(intermediate_reg_0[5660]),.o(intermediate_reg_1[2830]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5659]),.i2(intermediate_reg_0[5658]),.o(intermediate_reg_1[2829])); 
fsm fsm_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5657]),.i2(intermediate_reg_0[5656]),.o(intermediate_reg_1[2828])); 
fsm fsm_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5655]),.i2(intermediate_reg_0[5654]),.o(intermediate_reg_1[2827])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5653]),.i2(intermediate_reg_0[5652]),.o(intermediate_reg_1[2826]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5651]),.i2(intermediate_reg_0[5650]),.o(intermediate_reg_1[2825]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5649]),.i2(intermediate_reg_0[5648]),.o(intermediate_reg_1[2824])); 
fsm fsm_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5647]),.i2(intermediate_reg_0[5646]),.o(intermediate_reg_1[2823])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5645]),.i2(intermediate_reg_0[5644]),.o(intermediate_reg_1[2822])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5643]),.i2(intermediate_reg_0[5642]),.o(intermediate_reg_1[2821]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5641]),.i2(intermediate_reg_0[5640]),.o(intermediate_reg_1[2820])); 
fsm fsm_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5639]),.i2(intermediate_reg_0[5638]),.o(intermediate_reg_1[2819])); 
fsm fsm_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5637]),.i2(intermediate_reg_0[5636]),.o(intermediate_reg_1[2818])); 
fsm fsm_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5635]),.i2(intermediate_reg_0[5634]),.o(intermediate_reg_1[2817])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5633]),.i2(intermediate_reg_0[5632]),.o(intermediate_reg_1[2816]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5631]),.i2(intermediate_reg_0[5630]),.o(intermediate_reg_1[2815])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5629]),.i2(intermediate_reg_0[5628]),.o(intermediate_reg_1[2814]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5627]),.i2(intermediate_reg_0[5626]),.o(intermediate_reg_1[2813])); 
mux_module mux_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5625]),.i2(intermediate_reg_0[5624]),.o(intermediate_reg_1[2812]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5623]),.i2(intermediate_reg_0[5622]),.o(intermediate_reg_1[2811])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5621]),.i2(intermediate_reg_0[5620]),.o(intermediate_reg_1[2810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5619]),.i2(intermediate_reg_0[5618]),.o(intermediate_reg_1[2809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5617]),.i2(intermediate_reg_0[5616]),.o(intermediate_reg_1[2808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5615]),.i2(intermediate_reg_0[5614]),.o(intermediate_reg_1[2807]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5613]),.i2(intermediate_reg_0[5612]),.o(intermediate_reg_1[2806])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5611]),.i2(intermediate_reg_0[5610]),.o(intermediate_reg_1[2805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5609]),.i2(intermediate_reg_0[5608]),.o(intermediate_reg_1[2804]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5607]),.i2(intermediate_reg_0[5606]),.o(intermediate_reg_1[2803])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5605]),.i2(intermediate_reg_0[5604]),.o(intermediate_reg_1[2802])); 
fsm fsm_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5603]),.i2(intermediate_reg_0[5602]),.o(intermediate_reg_1[2801])); 
fsm fsm_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5601]),.i2(intermediate_reg_0[5600]),.o(intermediate_reg_1[2800])); 
mux_module mux_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5599]),.i2(intermediate_reg_0[5598]),.o(intermediate_reg_1[2799]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5597]),.i2(intermediate_reg_0[5596]),.o(intermediate_reg_1[2798]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5595]),.i2(intermediate_reg_0[5594]),.o(intermediate_reg_1[2797]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5593]),.i2(intermediate_reg_0[5592]),.o(intermediate_reg_1[2796]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5591]),.i2(intermediate_reg_0[5590]),.o(intermediate_reg_1[2795])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5589]),.i2(intermediate_reg_0[5588]),.o(intermediate_reg_1[2794])); 
fsm fsm_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5587]),.i2(intermediate_reg_0[5586]),.o(intermediate_reg_1[2793])); 
fsm fsm_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5585]),.i2(intermediate_reg_0[5584]),.o(intermediate_reg_1[2792])); 
fsm fsm_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5583]),.i2(intermediate_reg_0[5582]),.o(intermediate_reg_1[2791])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5581]),.i2(intermediate_reg_0[5580]),.o(intermediate_reg_1[2790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5579]),.i2(intermediate_reg_0[5578]),.o(intermediate_reg_1[2789]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5577]),.i2(intermediate_reg_0[5576]),.o(intermediate_reg_1[2788])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5575]),.i2(intermediate_reg_0[5574]),.o(intermediate_reg_1[2787]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5573]),.i2(intermediate_reg_0[5572]),.o(intermediate_reg_1[2786]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5571]),.i2(intermediate_reg_0[5570]),.o(intermediate_reg_1[2785]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5569]),.i2(intermediate_reg_0[5568]),.o(intermediate_reg_1[2784])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5567]),.i2(intermediate_reg_0[5566]),.o(intermediate_reg_1[2783]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5565]),.i2(intermediate_reg_0[5564]),.o(intermediate_reg_1[2782])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5563]),.i2(intermediate_reg_0[5562]),.o(intermediate_reg_1[2781])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5561]),.i2(intermediate_reg_0[5560]),.o(intermediate_reg_1[2780]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5559]),.i2(intermediate_reg_0[5558]),.o(intermediate_reg_1[2779]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5557]),.i2(intermediate_reg_0[5556]),.o(intermediate_reg_1[2778]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5555]),.i2(intermediate_reg_0[5554]),.o(intermediate_reg_1[2777])); 
fsm fsm_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5553]),.i2(intermediate_reg_0[5552]),.o(intermediate_reg_1[2776])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5551]),.i2(intermediate_reg_0[5550]),.o(intermediate_reg_1[2775]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5549]),.i2(intermediate_reg_0[5548]),.o(intermediate_reg_1[2774])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5547]),.i2(intermediate_reg_0[5546]),.o(intermediate_reg_1[2773]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5545]),.i2(intermediate_reg_0[5544]),.o(intermediate_reg_1[2772])); 
fsm fsm_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5543]),.i2(intermediate_reg_0[5542]),.o(intermediate_reg_1[2771])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5541]),.i2(intermediate_reg_0[5540]),.o(intermediate_reg_1[2770])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5539]),.i2(intermediate_reg_0[5538]),.o(intermediate_reg_1[2769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5537]),.i2(intermediate_reg_0[5536]),.o(intermediate_reg_1[2768]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5535]),.i2(intermediate_reg_0[5534]),.o(intermediate_reg_1[2767]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5533]),.i2(intermediate_reg_0[5532]),.o(intermediate_reg_1[2766])); 
fsm fsm_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5531]),.i2(intermediate_reg_0[5530]),.o(intermediate_reg_1[2765])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5529]),.i2(intermediate_reg_0[5528]),.o(intermediate_reg_1[2764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5527]),.i2(intermediate_reg_0[5526]),.o(intermediate_reg_1[2763]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5525]),.i2(intermediate_reg_0[5524]),.o(intermediate_reg_1[2762]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5523]),.i2(intermediate_reg_0[5522]),.o(intermediate_reg_1[2761])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5521]),.i2(intermediate_reg_0[5520]),.o(intermediate_reg_1[2760]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5519]),.i2(intermediate_reg_0[5518]),.o(intermediate_reg_1[2759])); 
fsm fsm_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5517]),.i2(intermediate_reg_0[5516]),.o(intermediate_reg_1[2758])); 
fsm fsm_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5515]),.i2(intermediate_reg_0[5514]),.o(intermediate_reg_1[2757])); 
mux_module mux_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5513]),.i2(intermediate_reg_0[5512]),.o(intermediate_reg_1[2756]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5511]),.i2(intermediate_reg_0[5510]),.o(intermediate_reg_1[2755])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5509]),.i2(intermediate_reg_0[5508]),.o(intermediate_reg_1[2754]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5507]),.i2(intermediate_reg_0[5506]),.o(intermediate_reg_1[2753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5505]),.i2(intermediate_reg_0[5504]),.o(intermediate_reg_1[2752]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5503]),.i2(intermediate_reg_0[5502]),.o(intermediate_reg_1[2751]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5501]),.i2(intermediate_reg_0[5500]),.o(intermediate_reg_1[2750])); 
mux_module mux_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5499]),.i2(intermediate_reg_0[5498]),.o(intermediate_reg_1[2749]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5497]),.i2(intermediate_reg_0[5496]),.o(intermediate_reg_1[2748]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5495]),.i2(intermediate_reg_0[5494]),.o(intermediate_reg_1[2747]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5493]),.i2(intermediate_reg_0[5492]),.o(intermediate_reg_1[2746])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5491]),.i2(intermediate_reg_0[5490]),.o(intermediate_reg_1[2745]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5489]),.i2(intermediate_reg_0[5488]),.o(intermediate_reg_1[2744])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5487]),.i2(intermediate_reg_0[5486]),.o(intermediate_reg_1[2743]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5485]),.i2(intermediate_reg_0[5484]),.o(intermediate_reg_1[2742]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5483]),.i2(intermediate_reg_0[5482]),.o(intermediate_reg_1[2741]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5481]),.i2(intermediate_reg_0[5480]),.o(intermediate_reg_1[2740])); 
fsm fsm_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5479]),.i2(intermediate_reg_0[5478]),.o(intermediate_reg_1[2739])); 
fsm fsm_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5477]),.i2(intermediate_reg_0[5476]),.o(intermediate_reg_1[2738])); 
fsm fsm_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5475]),.i2(intermediate_reg_0[5474]),.o(intermediate_reg_1[2737])); 
fsm fsm_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5473]),.i2(intermediate_reg_0[5472]),.o(intermediate_reg_1[2736])); 
mux_module mux_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5471]),.i2(intermediate_reg_0[5470]),.o(intermediate_reg_1[2735]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5469]),.i2(intermediate_reg_0[5468]),.o(intermediate_reg_1[2734])); 
fsm fsm_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5467]),.i2(intermediate_reg_0[5466]),.o(intermediate_reg_1[2733])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5465]),.i2(intermediate_reg_0[5464]),.o(intermediate_reg_1[2732]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5463]),.i2(intermediate_reg_0[5462]),.o(intermediate_reg_1[2731])); 
fsm fsm_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5461]),.i2(intermediate_reg_0[5460]),.o(intermediate_reg_1[2730])); 
mux_module mux_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5459]),.i2(intermediate_reg_0[5458]),.o(intermediate_reg_1[2729]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5457]),.i2(intermediate_reg_0[5456]),.o(intermediate_reg_1[2728])); 
mux_module mux_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5455]),.i2(intermediate_reg_0[5454]),.o(intermediate_reg_1[2727]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5453]),.i2(intermediate_reg_0[5452]),.o(intermediate_reg_1[2726])); 
fsm fsm_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5451]),.i2(intermediate_reg_0[5450]),.o(intermediate_reg_1[2725])); 
mux_module mux_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5449]),.i2(intermediate_reg_0[5448]),.o(intermediate_reg_1[2724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5447]),.i2(intermediate_reg_0[5446]),.o(intermediate_reg_1[2723]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5445]),.i2(intermediate_reg_0[5444]),.o(intermediate_reg_1[2722])); 
mux_module mux_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5443]),.i2(intermediate_reg_0[5442]),.o(intermediate_reg_1[2721]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5441]),.i2(intermediate_reg_0[5440]),.o(intermediate_reg_1[2720]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5439]),.i2(intermediate_reg_0[5438]),.o(intermediate_reg_1[2719]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5437]),.i2(intermediate_reg_0[5436]),.o(intermediate_reg_1[2718])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5435]),.i2(intermediate_reg_0[5434]),.o(intermediate_reg_1[2717])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5433]),.i2(intermediate_reg_0[5432]),.o(intermediate_reg_1[2716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5431]),.i2(intermediate_reg_0[5430]),.o(intermediate_reg_1[2715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5429]),.i2(intermediate_reg_0[5428]),.o(intermediate_reg_1[2714]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5427]),.i2(intermediate_reg_0[5426]),.o(intermediate_reg_1[2713]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5425]),.i2(intermediate_reg_0[5424]),.o(intermediate_reg_1[2712]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5423]),.i2(intermediate_reg_0[5422]),.o(intermediate_reg_1[2711]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5421]),.i2(intermediate_reg_0[5420]),.o(intermediate_reg_1[2710])); 
fsm fsm_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5419]),.i2(intermediate_reg_0[5418]),.o(intermediate_reg_1[2709])); 
fsm fsm_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5417]),.i2(intermediate_reg_0[5416]),.o(intermediate_reg_1[2708])); 
fsm fsm_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5415]),.i2(intermediate_reg_0[5414]),.o(intermediate_reg_1[2707])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5413]),.i2(intermediate_reg_0[5412]),.o(intermediate_reg_1[2706])); 
fsm fsm_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5411]),.i2(intermediate_reg_0[5410]),.o(intermediate_reg_1[2705])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5409]),.i2(intermediate_reg_0[5408]),.o(intermediate_reg_1[2704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5407]),.i2(intermediate_reg_0[5406]),.o(intermediate_reg_1[2703]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5405]),.i2(intermediate_reg_0[5404]),.o(intermediate_reg_1[2702])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5403]),.i2(intermediate_reg_0[5402]),.o(intermediate_reg_1[2701]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5401]),.i2(intermediate_reg_0[5400]),.o(intermediate_reg_1[2700])); 
fsm fsm_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5399]),.i2(intermediate_reg_0[5398]),.o(intermediate_reg_1[2699])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5397]),.i2(intermediate_reg_0[5396]),.o(intermediate_reg_1[2698]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5395]),.i2(intermediate_reg_0[5394]),.o(intermediate_reg_1[2697])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5393]),.i2(intermediate_reg_0[5392]),.o(intermediate_reg_1[2696]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5391]),.i2(intermediate_reg_0[5390]),.o(intermediate_reg_1[2695])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5389]),.i2(intermediate_reg_0[5388]),.o(intermediate_reg_1[2694])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5387]),.i2(intermediate_reg_0[5386]),.o(intermediate_reg_1[2693])); 
fsm fsm_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5385]),.i2(intermediate_reg_0[5384]),.o(intermediate_reg_1[2692])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5383]),.i2(intermediate_reg_0[5382]),.o(intermediate_reg_1[2691]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5381]),.i2(intermediate_reg_0[5380]),.o(intermediate_reg_1[2690])); 
mux_module mux_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5379]),.i2(intermediate_reg_0[5378]),.o(intermediate_reg_1[2689]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5377]),.i2(intermediate_reg_0[5376]),.o(intermediate_reg_1[2688])); 
fsm fsm_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5375]),.i2(intermediate_reg_0[5374]),.o(intermediate_reg_1[2687])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5373]),.i2(intermediate_reg_0[5372]),.o(intermediate_reg_1[2686]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5371]),.i2(intermediate_reg_0[5370]),.o(intermediate_reg_1[2685]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5369]),.i2(intermediate_reg_0[5368]),.o(intermediate_reg_1[2684])); 
mux_module mux_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5367]),.i2(intermediate_reg_0[5366]),.o(intermediate_reg_1[2683]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5365]),.i2(intermediate_reg_0[5364]),.o(intermediate_reg_1[2682])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5363]),.i2(intermediate_reg_0[5362]),.o(intermediate_reg_1[2681])); 
fsm fsm_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5361]),.i2(intermediate_reg_0[5360]),.o(intermediate_reg_1[2680])); 
fsm fsm_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5359]),.i2(intermediate_reg_0[5358]),.o(intermediate_reg_1[2679])); 
mux_module mux_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5357]),.i2(intermediate_reg_0[5356]),.o(intermediate_reg_1[2678]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5355]),.i2(intermediate_reg_0[5354]),.o(intermediate_reg_1[2677])); 
mux_module mux_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5353]),.i2(intermediate_reg_0[5352]),.o(intermediate_reg_1[2676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5351]),.i2(intermediate_reg_0[5350]),.o(intermediate_reg_1[2675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5349]),.i2(intermediate_reg_0[5348]),.o(intermediate_reg_1[2674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5347]),.i2(intermediate_reg_0[5346]),.o(intermediate_reg_1[2673]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5345]),.i2(intermediate_reg_0[5344]),.o(intermediate_reg_1[2672])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5343]),.i2(intermediate_reg_0[5342]),.o(intermediate_reg_1[2671]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5341]),.i2(intermediate_reg_0[5340]),.o(intermediate_reg_1[2670])); 
mux_module mux_module_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5339]),.i2(intermediate_reg_0[5338]),.o(intermediate_reg_1[2669]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5337]),.i2(intermediate_reg_0[5336]),.o(intermediate_reg_1[2668])); 
mux_module mux_module_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5335]),.i2(intermediate_reg_0[5334]),.o(intermediate_reg_1[2667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5333]),.i2(intermediate_reg_0[5332]),.o(intermediate_reg_1[2666]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5331]),.i2(intermediate_reg_0[5330]),.o(intermediate_reg_1[2665])); 
mux_module mux_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5329]),.i2(intermediate_reg_0[5328]),.o(intermediate_reg_1[2664]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5327]),.i2(intermediate_reg_0[5326]),.o(intermediate_reg_1[2663])); 
fsm fsm_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5325]),.i2(intermediate_reg_0[5324]),.o(intermediate_reg_1[2662])); 
mux_module mux_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5323]),.i2(intermediate_reg_0[5322]),.o(intermediate_reg_1[2661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5321]),.i2(intermediate_reg_0[5320]),.o(intermediate_reg_1[2660]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5319]),.i2(intermediate_reg_0[5318]),.o(intermediate_reg_1[2659])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5317]),.i2(intermediate_reg_0[5316]),.o(intermediate_reg_1[2658])); 
mux_module mux_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5315]),.i2(intermediate_reg_0[5314]),.o(intermediate_reg_1[2657]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5313]),.i2(intermediate_reg_0[5312]),.o(intermediate_reg_1[2656])); 
fsm fsm_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5311]),.i2(intermediate_reg_0[5310]),.o(intermediate_reg_1[2655])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5309]),.i2(intermediate_reg_0[5308]),.o(intermediate_reg_1[2654]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5307]),.i2(intermediate_reg_0[5306]),.o(intermediate_reg_1[2653])); 
fsm fsm_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5305]),.i2(intermediate_reg_0[5304]),.o(intermediate_reg_1[2652])); 
fsm fsm_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5303]),.i2(intermediate_reg_0[5302]),.o(intermediate_reg_1[2651])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5301]),.i2(intermediate_reg_0[5300]),.o(intermediate_reg_1[2650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5299]),.i2(intermediate_reg_0[5298]),.o(intermediate_reg_1[2649]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5297]),.i2(intermediate_reg_0[5296]),.o(intermediate_reg_1[2648])); 
fsm fsm_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5295]),.i2(intermediate_reg_0[5294]),.o(intermediate_reg_1[2647])); 
fsm fsm_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5293]),.i2(intermediate_reg_0[5292]),.o(intermediate_reg_1[2646])); 
fsm fsm_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5291]),.i2(intermediate_reg_0[5290]),.o(intermediate_reg_1[2645])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5289]),.i2(intermediate_reg_0[5288]),.o(intermediate_reg_1[2644])); 
fsm fsm_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5287]),.i2(intermediate_reg_0[5286]),.o(intermediate_reg_1[2643])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5285]),.i2(intermediate_reg_0[5284]),.o(intermediate_reg_1[2642])); 
mux_module mux_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5283]),.i2(intermediate_reg_0[5282]),.o(intermediate_reg_1[2641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5281]),.i2(intermediate_reg_0[5280]),.o(intermediate_reg_1[2640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5279]),.i2(intermediate_reg_0[5278]),.o(intermediate_reg_1[2639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5277]),.i2(intermediate_reg_0[5276]),.o(intermediate_reg_1[2638]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5275]),.i2(intermediate_reg_0[5274]),.o(intermediate_reg_1[2637]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5273]),.i2(intermediate_reg_0[5272]),.o(intermediate_reg_1[2636]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5271]),.i2(intermediate_reg_0[5270]),.o(intermediate_reg_1[2635])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5269]),.i2(intermediate_reg_0[5268]),.o(intermediate_reg_1[2634])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5267]),.i2(intermediate_reg_0[5266]),.o(intermediate_reg_1[2633])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5265]),.i2(intermediate_reg_0[5264]),.o(intermediate_reg_1[2632])); 
mux_module mux_module_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5263]),.i2(intermediate_reg_0[5262]),.o(intermediate_reg_1[2631]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5261]),.i2(intermediate_reg_0[5260]),.o(intermediate_reg_1[2630])); 
fsm fsm_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5259]),.i2(intermediate_reg_0[5258]),.o(intermediate_reg_1[2629])); 
mux_module mux_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5257]),.i2(intermediate_reg_0[5256]),.o(intermediate_reg_1[2628]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5255]),.i2(intermediate_reg_0[5254]),.o(intermediate_reg_1[2627]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5253]),.i2(intermediate_reg_0[5252]),.o(intermediate_reg_1[2626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5251]),.i2(intermediate_reg_0[5250]),.o(intermediate_reg_1[2625])); 
fsm fsm_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5249]),.i2(intermediate_reg_0[5248]),.o(intermediate_reg_1[2624])); 
fsm fsm_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5247]),.i2(intermediate_reg_0[5246]),.o(intermediate_reg_1[2623])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5245]),.i2(intermediate_reg_0[5244]),.o(intermediate_reg_1[2622])); 
mux_module mux_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5243]),.i2(intermediate_reg_0[5242]),.o(intermediate_reg_1[2621]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5241]),.i2(intermediate_reg_0[5240]),.o(intermediate_reg_1[2620])); 
fsm fsm_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5239]),.i2(intermediate_reg_0[5238]),.o(intermediate_reg_1[2619])); 
fsm fsm_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5237]),.i2(intermediate_reg_0[5236]),.o(intermediate_reg_1[2618])); 
fsm fsm_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5235]),.i2(intermediate_reg_0[5234]),.o(intermediate_reg_1[2617])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5233]),.i2(intermediate_reg_0[5232]),.o(intermediate_reg_1[2616])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5231]),.i2(intermediate_reg_0[5230]),.o(intermediate_reg_1[2615])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5229]),.i2(intermediate_reg_0[5228]),.o(intermediate_reg_1[2614])); 
mux_module mux_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5227]),.i2(intermediate_reg_0[5226]),.o(intermediate_reg_1[2613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5225]),.i2(intermediate_reg_0[5224]),.o(intermediate_reg_1[2612]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5223]),.i2(intermediate_reg_0[5222]),.o(intermediate_reg_1[2611]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5221]),.i2(intermediate_reg_0[5220]),.o(intermediate_reg_1[2610])); 
mux_module mux_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5219]),.i2(intermediate_reg_0[5218]),.o(intermediate_reg_1[2609]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5217]),.i2(intermediate_reg_0[5216]),.o(intermediate_reg_1[2608])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5215]),.i2(intermediate_reg_0[5214]),.o(intermediate_reg_1[2607]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5213]),.i2(intermediate_reg_0[5212]),.o(intermediate_reg_1[2606])); 
fsm fsm_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5211]),.i2(intermediate_reg_0[5210]),.o(intermediate_reg_1[2605])); 
mux_module mux_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5209]),.i2(intermediate_reg_0[5208]),.o(intermediate_reg_1[2604]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5207]),.i2(intermediate_reg_0[5206]),.o(intermediate_reg_1[2603])); 
fsm fsm_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5205]),.i2(intermediate_reg_0[5204]),.o(intermediate_reg_1[2602])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5203]),.i2(intermediate_reg_0[5202]),.o(intermediate_reg_1[2601]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5201]),.i2(intermediate_reg_0[5200]),.o(intermediate_reg_1[2600]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5199]),.i2(intermediate_reg_0[5198]),.o(intermediate_reg_1[2599])); 
mux_module mux_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5197]),.i2(intermediate_reg_0[5196]),.o(intermediate_reg_1[2598]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5195]),.i2(intermediate_reg_0[5194]),.o(intermediate_reg_1[2597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5193]),.i2(intermediate_reg_0[5192]),.o(intermediate_reg_1[2596]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5191]),.i2(intermediate_reg_0[5190]),.o(intermediate_reg_1[2595]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5189]),.i2(intermediate_reg_0[5188]),.o(intermediate_reg_1[2594])); 
fsm fsm_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5187]),.i2(intermediate_reg_0[5186]),.o(intermediate_reg_1[2593])); 
fsm fsm_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5185]),.i2(intermediate_reg_0[5184]),.o(intermediate_reg_1[2592])); 
mux_module mux_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5183]),.i2(intermediate_reg_0[5182]),.o(intermediate_reg_1[2591]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5181]),.i2(intermediate_reg_0[5180]),.o(intermediate_reg_1[2590]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5179]),.i2(intermediate_reg_0[5178]),.o(intermediate_reg_1[2589]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5177]),.i2(intermediate_reg_0[5176]),.o(intermediate_reg_1[2588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5175]),.i2(intermediate_reg_0[5174]),.o(intermediate_reg_1[2587]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5173]),.i2(intermediate_reg_0[5172]),.o(intermediate_reg_1[2586])); 
fsm fsm_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5171]),.i2(intermediate_reg_0[5170]),.o(intermediate_reg_1[2585])); 
fsm fsm_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5169]),.i2(intermediate_reg_0[5168]),.o(intermediate_reg_1[2584])); 
fsm fsm_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5167]),.i2(intermediate_reg_0[5166]),.o(intermediate_reg_1[2583])); 
fsm fsm_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5165]),.i2(intermediate_reg_0[5164]),.o(intermediate_reg_1[2582])); 
mux_module mux_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5163]),.i2(intermediate_reg_0[5162]),.o(intermediate_reg_1[2581]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5161]),.i2(intermediate_reg_0[5160]),.o(intermediate_reg_1[2580]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5159]),.i2(intermediate_reg_0[5158]),.o(intermediate_reg_1[2579])); 
fsm fsm_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5157]),.i2(intermediate_reg_0[5156]),.o(intermediate_reg_1[2578])); 
mux_module mux_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5155]),.i2(intermediate_reg_0[5154]),.o(intermediate_reg_1[2577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5153]),.i2(intermediate_reg_0[5152]),.o(intermediate_reg_1[2576]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5151]),.i2(intermediate_reg_0[5150]),.o(intermediate_reg_1[2575])); 
mux_module mux_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5149]),.i2(intermediate_reg_0[5148]),.o(intermediate_reg_1[2574]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5147]),.i2(intermediate_reg_0[5146]),.o(intermediate_reg_1[2573]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5145]),.i2(intermediate_reg_0[5144]),.o(intermediate_reg_1[2572])); 
mux_module mux_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5143]),.i2(intermediate_reg_0[5142]),.o(intermediate_reg_1[2571]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5141]),.i2(intermediate_reg_0[5140]),.o(intermediate_reg_1[2570])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5139]),.i2(intermediate_reg_0[5138]),.o(intermediate_reg_1[2569]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5137]),.i2(intermediate_reg_0[5136]),.o(intermediate_reg_1[2568])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5135]),.i2(intermediate_reg_0[5134]),.o(intermediate_reg_1[2567]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5133]),.i2(intermediate_reg_0[5132]),.o(intermediate_reg_1[2566])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5131]),.i2(intermediate_reg_0[5130]),.o(intermediate_reg_1[2565]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5129]),.i2(intermediate_reg_0[5128]),.o(intermediate_reg_1[2564])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5127]),.i2(intermediate_reg_0[5126]),.o(intermediate_reg_1[2563]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5125]),.i2(intermediate_reg_0[5124]),.o(intermediate_reg_1[2562]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5123]),.i2(intermediate_reg_0[5122]),.o(intermediate_reg_1[2561])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5121]),.i2(intermediate_reg_0[5120]),.o(intermediate_reg_1[2560])); 
fsm fsm_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5119]),.i2(intermediate_reg_0[5118]),.o(intermediate_reg_1[2559])); 
fsm fsm_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5117]),.i2(intermediate_reg_0[5116]),.o(intermediate_reg_1[2558])); 
fsm fsm_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5115]),.i2(intermediate_reg_0[5114]),.o(intermediate_reg_1[2557])); 
mux_module mux_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5113]),.i2(intermediate_reg_0[5112]),.o(intermediate_reg_1[2556]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5111]),.i2(intermediate_reg_0[5110]),.o(intermediate_reg_1[2555])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5109]),.i2(intermediate_reg_0[5108]),.o(intermediate_reg_1[2554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5107]),.i2(intermediate_reg_0[5106]),.o(intermediate_reg_1[2553]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5105]),.i2(intermediate_reg_0[5104]),.o(intermediate_reg_1[2552])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5103]),.i2(intermediate_reg_0[5102]),.o(intermediate_reg_1[2551]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5101]),.i2(intermediate_reg_0[5100]),.o(intermediate_reg_1[2550])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5099]),.i2(intermediate_reg_0[5098]),.o(intermediate_reg_1[2549]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5097]),.i2(intermediate_reg_0[5096]),.o(intermediate_reg_1[2548])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5095]),.i2(intermediate_reg_0[5094]),.o(intermediate_reg_1[2547]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5093]),.i2(intermediate_reg_0[5092]),.o(intermediate_reg_1[2546])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5091]),.i2(intermediate_reg_0[5090]),.o(intermediate_reg_1[2545]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5089]),.i2(intermediate_reg_0[5088]),.o(intermediate_reg_1[2544])); 
mux_module mux_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5087]),.i2(intermediate_reg_0[5086]),.o(intermediate_reg_1[2543]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5085]),.i2(intermediate_reg_0[5084]),.o(intermediate_reg_1[2542]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5083]),.i2(intermediate_reg_0[5082]),.o(intermediate_reg_1[2541]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5081]),.i2(intermediate_reg_0[5080]),.o(intermediate_reg_1[2540])); 
mux_module mux_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5079]),.i2(intermediate_reg_0[5078]),.o(intermediate_reg_1[2539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5077]),.i2(intermediate_reg_0[5076]),.o(intermediate_reg_1[2538]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5075]),.i2(intermediate_reg_0[5074]),.o(intermediate_reg_1[2537])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5073]),.i2(intermediate_reg_0[5072]),.o(intermediate_reg_1[2536])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5071]),.i2(intermediate_reg_0[5070]),.o(intermediate_reg_1[2535])); 
fsm fsm_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5069]),.i2(intermediate_reg_0[5068]),.o(intermediate_reg_1[2534])); 
mux_module mux_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5067]),.i2(intermediate_reg_0[5066]),.o(intermediate_reg_1[2533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5065]),.i2(intermediate_reg_0[5064]),.o(intermediate_reg_1[2532]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5063]),.i2(intermediate_reg_0[5062]),.o(intermediate_reg_1[2531])); 
fsm fsm_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5061]),.i2(intermediate_reg_0[5060]),.o(intermediate_reg_1[2530])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5059]),.i2(intermediate_reg_0[5058]),.o(intermediate_reg_1[2529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5057]),.i2(intermediate_reg_0[5056]),.o(intermediate_reg_1[2528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5055]),.i2(intermediate_reg_0[5054]),.o(intermediate_reg_1[2527]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5053]),.i2(intermediate_reg_0[5052]),.o(intermediate_reg_1[2526])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5051]),.i2(intermediate_reg_0[5050]),.o(intermediate_reg_1[2525]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5049]),.i2(intermediate_reg_0[5048]),.o(intermediate_reg_1[2524])); 
fsm fsm_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5047]),.i2(intermediate_reg_0[5046]),.o(intermediate_reg_1[2523])); 
mux_module mux_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5045]),.i2(intermediate_reg_0[5044]),.o(intermediate_reg_1[2522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5043]),.i2(intermediate_reg_0[5042]),.o(intermediate_reg_1[2521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5041]),.i2(intermediate_reg_0[5040]),.o(intermediate_reg_1[2520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5039]),.i2(intermediate_reg_0[5038]),.o(intermediate_reg_1[2519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5037]),.i2(intermediate_reg_0[5036]),.o(intermediate_reg_1[2518]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5035]),.i2(intermediate_reg_0[5034]),.o(intermediate_reg_1[2517]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5033]),.i2(intermediate_reg_0[5032]),.o(intermediate_reg_1[2516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5031]),.i2(intermediate_reg_0[5030]),.o(intermediate_reg_1[2515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5029]),.i2(intermediate_reg_0[5028]),.o(intermediate_reg_1[2514]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5027]),.i2(intermediate_reg_0[5026]),.o(intermediate_reg_1[2513]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5025]),.i2(intermediate_reg_0[5024]),.o(intermediate_reg_1[2512])); 
fsm fsm_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5023]),.i2(intermediate_reg_0[5022]),.o(intermediate_reg_1[2511])); 
mux_module mux_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5021]),.i2(intermediate_reg_0[5020]),.o(intermediate_reg_1[2510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5019]),.i2(intermediate_reg_0[5018]),.o(intermediate_reg_1[2509]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5017]),.i2(intermediate_reg_0[5016]),.o(intermediate_reg_1[2508])); 
fsm fsm_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5015]),.i2(intermediate_reg_0[5014]),.o(intermediate_reg_1[2507])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5013]),.i2(intermediate_reg_0[5012]),.o(intermediate_reg_1[2506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5011]),.i2(intermediate_reg_0[5010]),.o(intermediate_reg_1[2505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5009]),.i2(intermediate_reg_0[5008]),.o(intermediate_reg_1[2504]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5007]),.i2(intermediate_reg_0[5006]),.o(intermediate_reg_1[2503]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5005]),.i2(intermediate_reg_0[5004]),.o(intermediate_reg_1[2502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5003]),.i2(intermediate_reg_0[5002]),.o(intermediate_reg_1[2501]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5001]),.i2(intermediate_reg_0[5000]),.o(intermediate_reg_1[2500])); 
fsm fsm_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4999]),.i2(intermediate_reg_0[4998]),.o(intermediate_reg_1[2499])); 
mux_module mux_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4997]),.i2(intermediate_reg_0[4996]),.o(intermediate_reg_1[2498]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4995]),.i2(intermediate_reg_0[4994]),.o(intermediate_reg_1[2497])); 
fsm fsm_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4993]),.i2(intermediate_reg_0[4992]),.o(intermediate_reg_1[2496])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4991]),.i2(intermediate_reg_0[4990]),.o(intermediate_reg_1[2495]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4989]),.i2(intermediate_reg_0[4988]),.o(intermediate_reg_1[2494])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4987]),.i2(intermediate_reg_0[4986]),.o(intermediate_reg_1[2493])); 
mux_module mux_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4985]),.i2(intermediate_reg_0[4984]),.o(intermediate_reg_1[2492]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4983]),.i2(intermediate_reg_0[4982]),.o(intermediate_reg_1[2491])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4981]),.i2(intermediate_reg_0[4980]),.o(intermediate_reg_1[2490]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4979]),.i2(intermediate_reg_0[4978]),.o(intermediate_reg_1[2489])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4977]),.i2(intermediate_reg_0[4976]),.o(intermediate_reg_1[2488]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4975]),.i2(intermediate_reg_0[4974]),.o(intermediate_reg_1[2487])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4973]),.i2(intermediate_reg_0[4972]),.o(intermediate_reg_1[2486])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4971]),.i2(intermediate_reg_0[4970]),.o(intermediate_reg_1[2485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4969]),.i2(intermediate_reg_0[4968]),.o(intermediate_reg_1[2484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4967]),.i2(intermediate_reg_0[4966]),.o(intermediate_reg_1[2483]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4965]),.i2(intermediate_reg_0[4964]),.o(intermediate_reg_1[2482]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4963]),.i2(intermediate_reg_0[4962]),.o(intermediate_reg_1[2481])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4961]),.i2(intermediate_reg_0[4960]),.o(intermediate_reg_1[2480])); 
fsm fsm_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4959]),.i2(intermediate_reg_0[4958]),.o(intermediate_reg_1[2479])); 
fsm fsm_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4957]),.i2(intermediate_reg_0[4956]),.o(intermediate_reg_1[2478])); 
fsm fsm_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4955]),.i2(intermediate_reg_0[4954]),.o(intermediate_reg_1[2477])); 
fsm fsm_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4953]),.i2(intermediate_reg_0[4952]),.o(intermediate_reg_1[2476])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4951]),.i2(intermediate_reg_0[4950]),.o(intermediate_reg_1[2475]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4949]),.i2(intermediate_reg_0[4948]),.o(intermediate_reg_1[2474])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4947]),.i2(intermediate_reg_0[4946]),.o(intermediate_reg_1[2473]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4945]),.i2(intermediate_reg_0[4944]),.o(intermediate_reg_1[2472]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4943]),.i2(intermediate_reg_0[4942]),.o(intermediate_reg_1[2471]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4941]),.i2(intermediate_reg_0[4940]),.o(intermediate_reg_1[2470])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4939]),.i2(intermediate_reg_0[4938]),.o(intermediate_reg_1[2469]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4937]),.i2(intermediate_reg_0[4936]),.o(intermediate_reg_1[2468])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4935]),.i2(intermediate_reg_0[4934]),.o(intermediate_reg_1[2467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4933]),.i2(intermediate_reg_0[4932]),.o(intermediate_reg_1[2466]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4931]),.i2(intermediate_reg_0[4930]),.o(intermediate_reg_1[2465])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4929]),.i2(intermediate_reg_0[4928]),.o(intermediate_reg_1[2464])); 
fsm fsm_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4927]),.i2(intermediate_reg_0[4926]),.o(intermediate_reg_1[2463])); 
fsm fsm_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4925]),.i2(intermediate_reg_0[4924]),.o(intermediate_reg_1[2462])); 
mux_module mux_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4923]),.i2(intermediate_reg_0[4922]),.o(intermediate_reg_1[2461]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4921]),.i2(intermediate_reg_0[4920]),.o(intermediate_reg_1[2460])); 
mux_module mux_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4919]),.i2(intermediate_reg_0[4918]),.o(intermediate_reg_1[2459]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4917]),.i2(intermediate_reg_0[4916]),.o(intermediate_reg_1[2458])); 
fsm fsm_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4915]),.i2(intermediate_reg_0[4914]),.o(intermediate_reg_1[2457])); 
mux_module mux_module_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4913]),.i2(intermediate_reg_0[4912]),.o(intermediate_reg_1[2456]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4911]),.i2(intermediate_reg_0[4910]),.o(intermediate_reg_1[2455])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4909]),.i2(intermediate_reg_0[4908]),.o(intermediate_reg_1[2454])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4907]),.i2(intermediate_reg_0[4906]),.o(intermediate_reg_1[2453]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4905]),.i2(intermediate_reg_0[4904]),.o(intermediate_reg_1[2452])); 
fsm fsm_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4903]),.i2(intermediate_reg_0[4902]),.o(intermediate_reg_1[2451])); 
mux_module mux_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4901]),.i2(intermediate_reg_0[4900]),.o(intermediate_reg_1[2450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4899]),.i2(intermediate_reg_0[4898]),.o(intermediate_reg_1[2449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4897]),.i2(intermediate_reg_0[4896]),.o(intermediate_reg_1[2448])); 
fsm fsm_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4895]),.i2(intermediate_reg_0[4894]),.o(intermediate_reg_1[2447])); 
fsm fsm_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4893]),.i2(intermediate_reg_0[4892]),.o(intermediate_reg_1[2446])); 
mux_module mux_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4891]),.i2(intermediate_reg_0[4890]),.o(intermediate_reg_1[2445]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4889]),.i2(intermediate_reg_0[4888]),.o(intermediate_reg_1[2444])); 
fsm fsm_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4887]),.i2(intermediate_reg_0[4886]),.o(intermediate_reg_1[2443])); 
mux_module mux_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4885]),.i2(intermediate_reg_0[4884]),.o(intermediate_reg_1[2442]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4883]),.i2(intermediate_reg_0[4882]),.o(intermediate_reg_1[2441]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4881]),.i2(intermediate_reg_0[4880]),.o(intermediate_reg_1[2440])); 
fsm fsm_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4879]),.i2(intermediate_reg_0[4878]),.o(intermediate_reg_1[2439])); 
fsm fsm_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4877]),.i2(intermediate_reg_0[4876]),.o(intermediate_reg_1[2438])); 
fsm fsm_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4875]),.i2(intermediate_reg_0[4874]),.o(intermediate_reg_1[2437])); 
fsm fsm_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4873]),.i2(intermediate_reg_0[4872]),.o(intermediate_reg_1[2436])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4871]),.i2(intermediate_reg_0[4870]),.o(intermediate_reg_1[2435]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4869]),.i2(intermediate_reg_0[4868]),.o(intermediate_reg_1[2434]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4867]),.i2(intermediate_reg_0[4866]),.o(intermediate_reg_1[2433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4865]),.i2(intermediate_reg_0[4864]),.o(intermediate_reg_1[2432]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4863]),.i2(intermediate_reg_0[4862]),.o(intermediate_reg_1[2431]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4861]),.i2(intermediate_reg_0[4860]),.o(intermediate_reg_1[2430]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4859]),.i2(intermediate_reg_0[4858]),.o(intermediate_reg_1[2429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4857]),.i2(intermediate_reg_0[4856]),.o(intermediate_reg_1[2428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4855]),.i2(intermediate_reg_0[4854]),.o(intermediate_reg_1[2427]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4853]),.i2(intermediate_reg_0[4852]),.o(intermediate_reg_1[2426])); 
fsm fsm_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4851]),.i2(intermediate_reg_0[4850]),.o(intermediate_reg_1[2425])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4849]),.i2(intermediate_reg_0[4848]),.o(intermediate_reg_1[2424]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4847]),.i2(intermediate_reg_0[4846]),.o(intermediate_reg_1[2423])); 
fsm fsm_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4845]),.i2(intermediate_reg_0[4844]),.o(intermediate_reg_1[2422])); 
fsm fsm_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4843]),.i2(intermediate_reg_0[4842]),.o(intermediate_reg_1[2421])); 
mux_module mux_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4841]),.i2(intermediate_reg_0[4840]),.o(intermediate_reg_1[2420]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4839]),.i2(intermediate_reg_0[4838]),.o(intermediate_reg_1[2419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4837]),.i2(intermediate_reg_0[4836]),.o(intermediate_reg_1[2418]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4835]),.i2(intermediate_reg_0[4834]),.o(intermediate_reg_1[2417])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4833]),.i2(intermediate_reg_0[4832]),.o(intermediate_reg_1[2416]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4831]),.i2(intermediate_reg_0[4830]),.o(intermediate_reg_1[2415]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4829]),.i2(intermediate_reg_0[4828]),.o(intermediate_reg_1[2414]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4827]),.i2(intermediate_reg_0[4826]),.o(intermediate_reg_1[2413]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4825]),.i2(intermediate_reg_0[4824]),.o(intermediate_reg_1[2412]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4823]),.i2(intermediate_reg_0[4822]),.o(intermediate_reg_1[2411]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4821]),.i2(intermediate_reg_0[4820]),.o(intermediate_reg_1[2410]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4819]),.i2(intermediate_reg_0[4818]),.o(intermediate_reg_1[2409]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4817]),.i2(intermediate_reg_0[4816]),.o(intermediate_reg_1[2408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4815]),.i2(intermediate_reg_0[4814]),.o(intermediate_reg_1[2407]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4813]),.i2(intermediate_reg_0[4812]),.o(intermediate_reg_1[2406]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4811]),.i2(intermediate_reg_0[4810]),.o(intermediate_reg_1[2405])); 
mux_module mux_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4809]),.i2(intermediate_reg_0[4808]),.o(intermediate_reg_1[2404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4807]),.i2(intermediate_reg_0[4806]),.o(intermediate_reg_1[2403])); 
mux_module mux_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4805]),.i2(intermediate_reg_0[4804]),.o(intermediate_reg_1[2402]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4803]),.i2(intermediate_reg_0[4802]),.o(intermediate_reg_1[2401])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4801]),.i2(intermediate_reg_0[4800]),.o(intermediate_reg_1[2400])); 
mux_module mux_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4799]),.i2(intermediate_reg_0[4798]),.o(intermediate_reg_1[2399]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4797]),.i2(intermediate_reg_0[4796]),.o(intermediate_reg_1[2398]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4795]),.i2(intermediate_reg_0[4794]),.o(intermediate_reg_1[2397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4793]),.i2(intermediate_reg_0[4792]),.o(intermediate_reg_1[2396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4791]),.i2(intermediate_reg_0[4790]),.o(intermediate_reg_1[2395]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4789]),.i2(intermediate_reg_0[4788]),.o(intermediate_reg_1[2394])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4787]),.i2(intermediate_reg_0[4786]),.o(intermediate_reg_1[2393]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4785]),.i2(intermediate_reg_0[4784]),.o(intermediate_reg_1[2392])); 
fsm fsm_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4783]),.i2(intermediate_reg_0[4782]),.o(intermediate_reg_1[2391])); 
fsm fsm_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4781]),.i2(intermediate_reg_0[4780]),.o(intermediate_reg_1[2390])); 
mux_module mux_module_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4779]),.i2(intermediate_reg_0[4778]),.o(intermediate_reg_1[2389]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4777]),.i2(intermediate_reg_0[4776]),.o(intermediate_reg_1[2388])); 
mux_module mux_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4775]),.i2(intermediate_reg_0[4774]),.o(intermediate_reg_1[2387]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4773]),.i2(intermediate_reg_0[4772]),.o(intermediate_reg_1[2386]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4771]),.i2(intermediate_reg_0[4770]),.o(intermediate_reg_1[2385]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4769]),.i2(intermediate_reg_0[4768]),.o(intermediate_reg_1[2384]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4767]),.i2(intermediate_reg_0[4766]),.o(intermediate_reg_1[2383])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4765]),.i2(intermediate_reg_0[4764]),.o(intermediate_reg_1[2382]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4763]),.i2(intermediate_reg_0[4762]),.o(intermediate_reg_1[2381])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4761]),.i2(intermediate_reg_0[4760]),.o(intermediate_reg_1[2380])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4759]),.i2(intermediate_reg_0[4758]),.o(intermediate_reg_1[2379]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4757]),.i2(intermediate_reg_0[4756]),.o(intermediate_reg_1[2378])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4755]),.i2(intermediate_reg_0[4754]),.o(intermediate_reg_1[2377]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4753]),.i2(intermediate_reg_0[4752]),.o(intermediate_reg_1[2376]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4751]),.i2(intermediate_reg_0[4750]),.o(intermediate_reg_1[2375])); 
mux_module mux_module_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4749]),.i2(intermediate_reg_0[4748]),.o(intermediate_reg_1[2374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4747]),.i2(intermediate_reg_0[4746]),.o(intermediate_reg_1[2373]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4745]),.i2(intermediate_reg_0[4744]),.o(intermediate_reg_1[2372]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4743]),.i2(intermediate_reg_0[4742]),.o(intermediate_reg_1[2371])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4741]),.i2(intermediate_reg_0[4740]),.o(intermediate_reg_1[2370]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4739]),.i2(intermediate_reg_0[4738]),.o(intermediate_reg_1[2369]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4737]),.i2(intermediate_reg_0[4736]),.o(intermediate_reg_1[2368])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4735]),.i2(intermediate_reg_0[4734]),.o(intermediate_reg_1[2367]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4733]),.i2(intermediate_reg_0[4732]),.o(intermediate_reg_1[2366]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4731]),.i2(intermediate_reg_0[4730]),.o(intermediate_reg_1[2365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4729]),.i2(intermediate_reg_0[4728]),.o(intermediate_reg_1[2364]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4727]),.i2(intermediate_reg_0[4726]),.o(intermediate_reg_1[2363])); 
fsm fsm_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4725]),.i2(intermediate_reg_0[4724]),.o(intermediate_reg_1[2362])); 
fsm fsm_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4723]),.i2(intermediate_reg_0[4722]),.o(intermediate_reg_1[2361])); 
mux_module mux_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4721]),.i2(intermediate_reg_0[4720]),.o(intermediate_reg_1[2360]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4719]),.i2(intermediate_reg_0[4718]),.o(intermediate_reg_1[2359])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4717]),.i2(intermediate_reg_0[4716]),.o(intermediate_reg_1[2358])); 
mux_module mux_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4715]),.i2(intermediate_reg_0[4714]),.o(intermediate_reg_1[2357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4713]),.i2(intermediate_reg_0[4712]),.o(intermediate_reg_1[2356]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4711]),.i2(intermediate_reg_0[4710]),.o(intermediate_reg_1[2355])); 
mux_module mux_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4709]),.i2(intermediate_reg_0[4708]),.o(intermediate_reg_1[2354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4707]),.i2(intermediate_reg_0[4706]),.o(intermediate_reg_1[2353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4705]),.i2(intermediate_reg_0[4704]),.o(intermediate_reg_1[2352]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4703]),.i2(intermediate_reg_0[4702]),.o(intermediate_reg_1[2351])); 
mux_module mux_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4701]),.i2(intermediate_reg_0[4700]),.o(intermediate_reg_1[2350]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4699]),.i2(intermediate_reg_0[4698]),.o(intermediate_reg_1[2349]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4697]),.i2(intermediate_reg_0[4696]),.o(intermediate_reg_1[2348]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4695]),.i2(intermediate_reg_0[4694]),.o(intermediate_reg_1[2347]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4693]),.i2(intermediate_reg_0[4692]),.o(intermediate_reg_1[2346])); 
mux_module mux_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4691]),.i2(intermediate_reg_0[4690]),.o(intermediate_reg_1[2345]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4689]),.i2(intermediate_reg_0[4688]),.o(intermediate_reg_1[2344])); 
fsm fsm_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4687]),.i2(intermediate_reg_0[4686]),.o(intermediate_reg_1[2343])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4685]),.i2(intermediate_reg_0[4684]),.o(intermediate_reg_1[2342]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4683]),.i2(intermediate_reg_0[4682]),.o(intermediate_reg_1[2341])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4681]),.i2(intermediate_reg_0[4680]),.o(intermediate_reg_1[2340]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4679]),.i2(intermediate_reg_0[4678]),.o(intermediate_reg_1[2339])); 
mux_module mux_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4677]),.i2(intermediate_reg_0[4676]),.o(intermediate_reg_1[2338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4675]),.i2(intermediate_reg_0[4674]),.o(intermediate_reg_1[2337]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4673]),.i2(intermediate_reg_0[4672]),.o(intermediate_reg_1[2336])); 
fsm fsm_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4671]),.i2(intermediate_reg_0[4670]),.o(intermediate_reg_1[2335])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4669]),.i2(intermediate_reg_0[4668]),.o(intermediate_reg_1[2334]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4667]),.i2(intermediate_reg_0[4666]),.o(intermediate_reg_1[2333])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4665]),.i2(intermediate_reg_0[4664]),.o(intermediate_reg_1[2332]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4663]),.i2(intermediate_reg_0[4662]),.o(intermediate_reg_1[2331])); 
mux_module mux_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4661]),.i2(intermediate_reg_0[4660]),.o(intermediate_reg_1[2330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4659]),.i2(intermediate_reg_0[4658]),.o(intermediate_reg_1[2329]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4657]),.i2(intermediate_reg_0[4656]),.o(intermediate_reg_1[2328])); 
fsm fsm_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4655]),.i2(intermediate_reg_0[4654]),.o(intermediate_reg_1[2327])); 
fsm fsm_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4653]),.i2(intermediate_reg_0[4652]),.o(intermediate_reg_1[2326])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4651]),.i2(intermediate_reg_0[4650]),.o(intermediate_reg_1[2325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4649]),.i2(intermediate_reg_0[4648]),.o(intermediate_reg_1[2324]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4647]),.i2(intermediate_reg_0[4646]),.o(intermediate_reg_1[2323])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4645]),.i2(intermediate_reg_0[4644]),.o(intermediate_reg_1[2322])); 
fsm fsm_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4643]),.i2(intermediate_reg_0[4642]),.o(intermediate_reg_1[2321])); 
fsm fsm_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4641]),.i2(intermediate_reg_0[4640]),.o(intermediate_reg_1[2320])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4639]),.i2(intermediate_reg_0[4638]),.o(intermediate_reg_1[2319]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4637]),.i2(intermediate_reg_0[4636]),.o(intermediate_reg_1[2318])); 
fsm fsm_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4635]),.i2(intermediate_reg_0[4634]),.o(intermediate_reg_1[2317])); 
mux_module mux_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4633]),.i2(intermediate_reg_0[4632]),.o(intermediate_reg_1[2316]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4631]),.i2(intermediate_reg_0[4630]),.o(intermediate_reg_1[2315])); 
fsm fsm_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4629]),.i2(intermediate_reg_0[4628]),.o(intermediate_reg_1[2314])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4627]),.i2(intermediate_reg_0[4626]),.o(intermediate_reg_1[2313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4625]),.i2(intermediate_reg_0[4624]),.o(intermediate_reg_1[2312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4623]),.i2(intermediate_reg_0[4622]),.o(intermediate_reg_1[2311]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4621]),.i2(intermediate_reg_0[4620]),.o(intermediate_reg_1[2310])); 
fsm fsm_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4619]),.i2(intermediate_reg_0[4618]),.o(intermediate_reg_1[2309])); 
mux_module mux_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4617]),.i2(intermediate_reg_0[4616]),.o(intermediate_reg_1[2308]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4615]),.i2(intermediate_reg_0[4614]),.o(intermediate_reg_1[2307])); 
fsm fsm_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4613]),.i2(intermediate_reg_0[4612]),.o(intermediate_reg_1[2306])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4611]),.i2(intermediate_reg_0[4610]),.o(intermediate_reg_1[2305])); 
fsm fsm_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4609]),.i2(intermediate_reg_0[4608]),.o(intermediate_reg_1[2304])); 
fsm fsm_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4607]),.i2(intermediate_reg_0[4606]),.o(intermediate_reg_1[2303])); 
fsm fsm_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4605]),.i2(intermediate_reg_0[4604]),.o(intermediate_reg_1[2302])); 
fsm fsm_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4603]),.i2(intermediate_reg_0[4602]),.o(intermediate_reg_1[2301])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4601]),.i2(intermediate_reg_0[4600]),.o(intermediate_reg_1[2300])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4599]),.i2(intermediate_reg_0[4598]),.o(intermediate_reg_1[2299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4597]),.i2(intermediate_reg_0[4596]),.o(intermediate_reg_1[2298]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4595]),.i2(intermediate_reg_0[4594]),.o(intermediate_reg_1[2297])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4593]),.i2(intermediate_reg_0[4592]),.o(intermediate_reg_1[2296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4591]),.i2(intermediate_reg_0[4590]),.o(intermediate_reg_1[2295]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4589]),.i2(intermediate_reg_0[4588]),.o(intermediate_reg_1[2294]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4587]),.i2(intermediate_reg_0[4586]),.o(intermediate_reg_1[2293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4585]),.i2(intermediate_reg_0[4584]),.o(intermediate_reg_1[2292]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4583]),.i2(intermediate_reg_0[4582]),.o(intermediate_reg_1[2291])); 
mux_module mux_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4581]),.i2(intermediate_reg_0[4580]),.o(intermediate_reg_1[2290]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4579]),.i2(intermediate_reg_0[4578]),.o(intermediate_reg_1[2289])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4577]),.i2(intermediate_reg_0[4576]),.o(intermediate_reg_1[2288]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4575]),.i2(intermediate_reg_0[4574]),.o(intermediate_reg_1[2287])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4573]),.i2(intermediate_reg_0[4572]),.o(intermediate_reg_1[2286]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4571]),.i2(intermediate_reg_0[4570]),.o(intermediate_reg_1[2285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4569]),.i2(intermediate_reg_0[4568]),.o(intermediate_reg_1[2284]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4567]),.i2(intermediate_reg_0[4566]),.o(intermediate_reg_1[2283])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4565]),.i2(intermediate_reg_0[4564]),.o(intermediate_reg_1[2282])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4563]),.i2(intermediate_reg_0[4562]),.o(intermediate_reg_1[2281]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4561]),.i2(intermediate_reg_0[4560]),.o(intermediate_reg_1[2280])); 
fsm fsm_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4559]),.i2(intermediate_reg_0[4558]),.o(intermediate_reg_1[2279])); 
fsm fsm_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4557]),.i2(intermediate_reg_0[4556]),.o(intermediate_reg_1[2278])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4555]),.i2(intermediate_reg_0[4554]),.o(intermediate_reg_1[2277])); 
mux_module mux_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4553]),.i2(intermediate_reg_0[4552]),.o(intermediate_reg_1[2276]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4551]),.i2(intermediate_reg_0[4550]),.o(intermediate_reg_1[2275])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4549]),.i2(intermediate_reg_0[4548]),.o(intermediate_reg_1[2274]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4547]),.i2(intermediate_reg_0[4546]),.o(intermediate_reg_1[2273])); 
fsm fsm_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4545]),.i2(intermediate_reg_0[4544]),.o(intermediate_reg_1[2272])); 
fsm fsm_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4543]),.i2(intermediate_reg_0[4542]),.o(intermediate_reg_1[2271])); 
fsm fsm_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4541]),.i2(intermediate_reg_0[4540]),.o(intermediate_reg_1[2270])); 
fsm fsm_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4539]),.i2(intermediate_reg_0[4538]),.o(intermediate_reg_1[2269])); 
fsm fsm_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4537]),.i2(intermediate_reg_0[4536]),.o(intermediate_reg_1[2268])); 
mux_module mux_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4535]),.i2(intermediate_reg_0[4534]),.o(intermediate_reg_1[2267]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4533]),.i2(intermediate_reg_0[4532]),.o(intermediate_reg_1[2266]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4531]),.i2(intermediate_reg_0[4530]),.o(intermediate_reg_1[2265])); 
mux_module mux_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4529]),.i2(intermediate_reg_0[4528]),.o(intermediate_reg_1[2264]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4527]),.i2(intermediate_reg_0[4526]),.o(intermediate_reg_1[2263])); 
mux_module mux_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4525]),.i2(intermediate_reg_0[4524]),.o(intermediate_reg_1[2262]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4523]),.i2(intermediate_reg_0[4522]),.o(intermediate_reg_1[2261])); 
mux_module mux_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4521]),.i2(intermediate_reg_0[4520]),.o(intermediate_reg_1[2260]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4519]),.i2(intermediate_reg_0[4518]),.o(intermediate_reg_1[2259])); 
mux_module mux_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4517]),.i2(intermediate_reg_0[4516]),.o(intermediate_reg_1[2258]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4515]),.i2(intermediate_reg_0[4514]),.o(intermediate_reg_1[2257])); 
fsm fsm_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4513]),.i2(intermediate_reg_0[4512]),.o(intermediate_reg_1[2256])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4511]),.i2(intermediate_reg_0[4510]),.o(intermediate_reg_1[2255])); 
mux_module mux_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4509]),.i2(intermediate_reg_0[4508]),.o(intermediate_reg_1[2254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4507]),.i2(intermediate_reg_0[4506]),.o(intermediate_reg_1[2253]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4505]),.i2(intermediate_reg_0[4504]),.o(intermediate_reg_1[2252]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4503]),.i2(intermediate_reg_0[4502]),.o(intermediate_reg_1[2251])); 
mux_module mux_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4501]),.i2(intermediate_reg_0[4500]),.o(intermediate_reg_1[2250]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4499]),.i2(intermediate_reg_0[4498]),.o(intermediate_reg_1[2249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4497]),.i2(intermediate_reg_0[4496]),.o(intermediate_reg_1[2248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4495]),.i2(intermediate_reg_0[4494]),.o(intermediate_reg_1[2247]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4493]),.i2(intermediate_reg_0[4492]),.o(intermediate_reg_1[2246])); 
fsm fsm_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4491]),.i2(intermediate_reg_0[4490]),.o(intermediate_reg_1[2245])); 
fsm fsm_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4489]),.i2(intermediate_reg_0[4488]),.o(intermediate_reg_1[2244])); 
mux_module mux_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4487]),.i2(intermediate_reg_0[4486]),.o(intermediate_reg_1[2243]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4485]),.i2(intermediate_reg_0[4484]),.o(intermediate_reg_1[2242])); 
fsm fsm_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4483]),.i2(intermediate_reg_0[4482]),.o(intermediate_reg_1[2241])); 
fsm fsm_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4481]),.i2(intermediate_reg_0[4480]),.o(intermediate_reg_1[2240])); 
fsm fsm_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4479]),.i2(intermediate_reg_0[4478]),.o(intermediate_reg_1[2239])); 
fsm fsm_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4477]),.i2(intermediate_reg_0[4476]),.o(intermediate_reg_1[2238])); 
mux_module mux_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4475]),.i2(intermediate_reg_0[4474]),.o(intermediate_reg_1[2237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4473]),.i2(intermediate_reg_0[4472]),.o(intermediate_reg_1[2236]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4471]),.i2(intermediate_reg_0[4470]),.o(intermediate_reg_1[2235])); 
fsm fsm_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4469]),.i2(intermediate_reg_0[4468]),.o(intermediate_reg_1[2234])); 
mux_module mux_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4467]),.i2(intermediate_reg_0[4466]),.o(intermediate_reg_1[2233]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4465]),.i2(intermediate_reg_0[4464]),.o(intermediate_reg_1[2232])); 
fsm fsm_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4463]),.i2(intermediate_reg_0[4462]),.o(intermediate_reg_1[2231])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4461]),.i2(intermediate_reg_0[4460]),.o(intermediate_reg_1[2230]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4459]),.i2(intermediate_reg_0[4458]),.o(intermediate_reg_1[2229])); 
mux_module mux_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4457]),.i2(intermediate_reg_0[4456]),.o(intermediate_reg_1[2228]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4455]),.i2(intermediate_reg_0[4454]),.o(intermediate_reg_1[2227])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4453]),.i2(intermediate_reg_0[4452]),.o(intermediate_reg_1[2226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4451]),.i2(intermediate_reg_0[4450]),.o(intermediate_reg_1[2225]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4449]),.i2(intermediate_reg_0[4448]),.o(intermediate_reg_1[2224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4447]),.i2(intermediate_reg_0[4446]),.o(intermediate_reg_1[2223]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4445]),.i2(intermediate_reg_0[4444]),.o(intermediate_reg_1[2222]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4443]),.i2(intermediate_reg_0[4442]),.o(intermediate_reg_1[2221])); 
mux_module mux_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4441]),.i2(intermediate_reg_0[4440]),.o(intermediate_reg_1[2220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4439]),.i2(intermediate_reg_0[4438]),.o(intermediate_reg_1[2219]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4437]),.i2(intermediate_reg_0[4436]),.o(intermediate_reg_1[2218])); 
mux_module mux_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4435]),.i2(intermediate_reg_0[4434]),.o(intermediate_reg_1[2217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4433]),.i2(intermediate_reg_0[4432]),.o(intermediate_reg_1[2216]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4431]),.i2(intermediate_reg_0[4430]),.o(intermediate_reg_1[2215])); 
fsm fsm_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4429]),.i2(intermediate_reg_0[4428]),.o(intermediate_reg_1[2214])); 
fsm fsm_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4427]),.i2(intermediate_reg_0[4426]),.o(intermediate_reg_1[2213])); 
fsm fsm_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4425]),.i2(intermediate_reg_0[4424]),.o(intermediate_reg_1[2212])); 
fsm fsm_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4423]),.i2(intermediate_reg_0[4422]),.o(intermediate_reg_1[2211])); 
mux_module mux_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4421]),.i2(intermediate_reg_0[4420]),.o(intermediate_reg_1[2210]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4419]),.i2(intermediate_reg_0[4418]),.o(intermediate_reg_1[2209])); 
fsm fsm_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4417]),.i2(intermediate_reg_0[4416]),.o(intermediate_reg_1[2208])); 
fsm fsm_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4415]),.i2(intermediate_reg_0[4414]),.o(intermediate_reg_1[2207])); 
fsm fsm_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4413]),.i2(intermediate_reg_0[4412]),.o(intermediate_reg_1[2206])); 
fsm fsm_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4411]),.i2(intermediate_reg_0[4410]),.o(intermediate_reg_1[2205])); 
fsm fsm_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4409]),.i2(intermediate_reg_0[4408]),.o(intermediate_reg_1[2204])); 
fsm fsm_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4407]),.i2(intermediate_reg_0[4406]),.o(intermediate_reg_1[2203])); 
mux_module mux_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4405]),.i2(intermediate_reg_0[4404]),.o(intermediate_reg_1[2202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4403]),.i2(intermediate_reg_0[4402]),.o(intermediate_reg_1[2201]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4401]),.i2(intermediate_reg_0[4400]),.o(intermediate_reg_1[2200])); 
fsm fsm_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4399]),.i2(intermediate_reg_0[4398]),.o(intermediate_reg_1[2199])); 
mux_module mux_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4397]),.i2(intermediate_reg_0[4396]),.o(intermediate_reg_1[2198]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4395]),.i2(intermediate_reg_0[4394]),.o(intermediate_reg_1[2197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4393]),.i2(intermediate_reg_0[4392]),.o(intermediate_reg_1[2196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4391]),.i2(intermediate_reg_0[4390]),.o(intermediate_reg_1[2195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4389]),.i2(intermediate_reg_0[4388]),.o(intermediate_reg_1[2194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4387]),.i2(intermediate_reg_0[4386]),.o(intermediate_reg_1[2193]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4385]),.i2(intermediate_reg_0[4384]),.o(intermediate_reg_1[2192])); 
fsm fsm_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4383]),.i2(intermediate_reg_0[4382]),.o(intermediate_reg_1[2191])); 
fsm fsm_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4381]),.i2(intermediate_reg_0[4380]),.o(intermediate_reg_1[2190])); 
mux_module mux_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4379]),.i2(intermediate_reg_0[4378]),.o(intermediate_reg_1[2189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4377]),.i2(intermediate_reg_0[4376]),.o(intermediate_reg_1[2188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4375]),.i2(intermediate_reg_0[4374]),.o(intermediate_reg_1[2187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4373]),.i2(intermediate_reg_0[4372]),.o(intermediate_reg_1[2186]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4371]),.i2(intermediate_reg_0[4370]),.o(intermediate_reg_1[2185])); 
fsm fsm_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4369]),.i2(intermediate_reg_0[4368]),.o(intermediate_reg_1[2184])); 
fsm fsm_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4367]),.i2(intermediate_reg_0[4366]),.o(intermediate_reg_1[2183])); 
fsm fsm_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4365]),.i2(intermediate_reg_0[4364]),.o(intermediate_reg_1[2182])); 
fsm fsm_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4363]),.i2(intermediate_reg_0[4362]),.o(intermediate_reg_1[2181])); 
mux_module mux_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4361]),.i2(intermediate_reg_0[4360]),.o(intermediate_reg_1[2180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4359]),.i2(intermediate_reg_0[4358]),.o(intermediate_reg_1[2179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4357]),.i2(intermediate_reg_0[4356]),.o(intermediate_reg_1[2178]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4355]),.i2(intermediate_reg_0[4354]),.o(intermediate_reg_1[2177])); 
mux_module mux_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4353]),.i2(intermediate_reg_0[4352]),.o(intermediate_reg_1[2176]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4351]),.i2(intermediate_reg_0[4350]),.o(intermediate_reg_1[2175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4349]),.i2(intermediate_reg_0[4348]),.o(intermediate_reg_1[2174]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4347]),.i2(intermediate_reg_0[4346]),.o(intermediate_reg_1[2173])); 
fsm fsm_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4345]),.i2(intermediate_reg_0[4344]),.o(intermediate_reg_1[2172])); 
fsm fsm_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4343]),.i2(intermediate_reg_0[4342]),.o(intermediate_reg_1[2171])); 
fsm fsm_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4341]),.i2(intermediate_reg_0[4340]),.o(intermediate_reg_1[2170])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4339]),.i2(intermediate_reg_0[4338]),.o(intermediate_reg_1[2169])); 
fsm fsm_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4337]),.i2(intermediate_reg_0[4336]),.o(intermediate_reg_1[2168])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4335]),.i2(intermediate_reg_0[4334]),.o(intermediate_reg_1[2167]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4333]),.i2(intermediate_reg_0[4332]),.o(intermediate_reg_1[2166]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4331]),.i2(intermediate_reg_0[4330]),.o(intermediate_reg_1[2165])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4329]),.i2(intermediate_reg_0[4328]),.o(intermediate_reg_1[2164])); 
fsm fsm_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4327]),.i2(intermediate_reg_0[4326]),.o(intermediate_reg_1[2163])); 
mux_module mux_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4325]),.i2(intermediate_reg_0[4324]),.o(intermediate_reg_1[2162]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4323]),.i2(intermediate_reg_0[4322]),.o(intermediate_reg_1[2161])); 
fsm fsm_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4321]),.i2(intermediate_reg_0[4320]),.o(intermediate_reg_1[2160])); 
fsm fsm_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4319]),.i2(intermediate_reg_0[4318]),.o(intermediate_reg_1[2159])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4317]),.i2(intermediate_reg_0[4316]),.o(intermediate_reg_1[2158])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4315]),.i2(intermediate_reg_0[4314]),.o(intermediate_reg_1[2157]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4313]),.i2(intermediate_reg_0[4312]),.o(intermediate_reg_1[2156]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4311]),.i2(intermediate_reg_0[4310]),.o(intermediate_reg_1[2155]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4309]),.i2(intermediate_reg_0[4308]),.o(intermediate_reg_1[2154])); 
mux_module mux_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4307]),.i2(intermediate_reg_0[4306]),.o(intermediate_reg_1[2153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4305]),.i2(intermediate_reg_0[4304]),.o(intermediate_reg_1[2152]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4303]),.i2(intermediate_reg_0[4302]),.o(intermediate_reg_1[2151])); 
mux_module mux_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4301]),.i2(intermediate_reg_0[4300]),.o(intermediate_reg_1[2150]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4299]),.i2(intermediate_reg_0[4298]),.o(intermediate_reg_1[2149])); 
fsm fsm_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4297]),.i2(intermediate_reg_0[4296]),.o(intermediate_reg_1[2148])); 
fsm fsm_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4295]),.i2(intermediate_reg_0[4294]),.o(intermediate_reg_1[2147])); 
fsm fsm_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4293]),.i2(intermediate_reg_0[4292]),.o(intermediate_reg_1[2146])); 
fsm fsm_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4291]),.i2(intermediate_reg_0[4290]),.o(intermediate_reg_1[2145])); 
mux_module mux_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4289]),.i2(intermediate_reg_0[4288]),.o(intermediate_reg_1[2144]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4287]),.i2(intermediate_reg_0[4286]),.o(intermediate_reg_1[2143]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4285]),.i2(intermediate_reg_0[4284]),.o(intermediate_reg_1[2142])); 
mux_module mux_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4283]),.i2(intermediate_reg_0[4282]),.o(intermediate_reg_1[2141]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4281]),.i2(intermediate_reg_0[4280]),.o(intermediate_reg_1[2140]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4279]),.i2(intermediate_reg_0[4278]),.o(intermediate_reg_1[2139]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4277]),.i2(intermediate_reg_0[4276]),.o(intermediate_reg_1[2138])); 
mux_module mux_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4275]),.i2(intermediate_reg_0[4274]),.o(intermediate_reg_1[2137]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4273]),.i2(intermediate_reg_0[4272]),.o(intermediate_reg_1[2136])); 
mux_module mux_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4271]),.i2(intermediate_reg_0[4270]),.o(intermediate_reg_1[2135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4269]),.i2(intermediate_reg_0[4268]),.o(intermediate_reg_1[2134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4267]),.i2(intermediate_reg_0[4266]),.o(intermediate_reg_1[2133]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4265]),.i2(intermediate_reg_0[4264]),.o(intermediate_reg_1[2132])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4263]),.i2(intermediate_reg_0[4262]),.o(intermediate_reg_1[2131]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4261]),.i2(intermediate_reg_0[4260]),.o(intermediate_reg_1[2130])); 
fsm fsm_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4259]),.i2(intermediate_reg_0[4258]),.o(intermediate_reg_1[2129])); 
mux_module mux_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4257]),.i2(intermediate_reg_0[4256]),.o(intermediate_reg_1[2128]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4255]),.i2(intermediate_reg_0[4254]),.o(intermediate_reg_1[2127])); 
fsm fsm_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4253]),.i2(intermediate_reg_0[4252]),.o(intermediate_reg_1[2126])); 
mux_module mux_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4251]),.i2(intermediate_reg_0[4250]),.o(intermediate_reg_1[2125]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4249]),.i2(intermediate_reg_0[4248]),.o(intermediate_reg_1[2124]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4247]),.i2(intermediate_reg_0[4246]),.o(intermediate_reg_1[2123])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4245]),.i2(intermediate_reg_0[4244]),.o(intermediate_reg_1[2122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4243]),.i2(intermediate_reg_0[4242]),.o(intermediate_reg_1[2121]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4241]),.i2(intermediate_reg_0[4240]),.o(intermediate_reg_1[2120])); 
mux_module mux_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4239]),.i2(intermediate_reg_0[4238]),.o(intermediate_reg_1[2119]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4237]),.i2(intermediate_reg_0[4236]),.o(intermediate_reg_1[2118])); 
fsm fsm_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4235]),.i2(intermediate_reg_0[4234]),.o(intermediate_reg_1[2117])); 
fsm fsm_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4233]),.i2(intermediate_reg_0[4232]),.o(intermediate_reg_1[2116])); 
mux_module mux_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4231]),.i2(intermediate_reg_0[4230]),.o(intermediate_reg_1[2115]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4229]),.i2(intermediate_reg_0[4228]),.o(intermediate_reg_1[2114]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4227]),.i2(intermediate_reg_0[4226]),.o(intermediate_reg_1[2113])); 
mux_module mux_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4225]),.i2(intermediate_reg_0[4224]),.o(intermediate_reg_1[2112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4223]),.i2(intermediate_reg_0[4222]),.o(intermediate_reg_1[2111]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4221]),.i2(intermediate_reg_0[4220]),.o(intermediate_reg_1[2110]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4219]),.i2(intermediate_reg_0[4218]),.o(intermediate_reg_1[2109])); 
fsm fsm_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4217]),.i2(intermediate_reg_0[4216]),.o(intermediate_reg_1[2108])); 
mux_module mux_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4215]),.i2(intermediate_reg_0[4214]),.o(intermediate_reg_1[2107]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4213]),.i2(intermediate_reg_0[4212]),.o(intermediate_reg_1[2106])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4211]),.i2(intermediate_reg_0[4210]),.o(intermediate_reg_1[2105]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4209]),.i2(intermediate_reg_0[4208]),.o(intermediate_reg_1[2104])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4207]),.i2(intermediate_reg_0[4206]),.o(intermediate_reg_1[2103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4205]),.i2(intermediate_reg_0[4204]),.o(intermediate_reg_1[2102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4203]),.i2(intermediate_reg_0[4202]),.o(intermediate_reg_1[2101]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4201]),.i2(intermediate_reg_0[4200]),.o(intermediate_reg_1[2100])); 
mux_module mux_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4199]),.i2(intermediate_reg_0[4198]),.o(intermediate_reg_1[2099]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4197]),.i2(intermediate_reg_0[4196]),.o(intermediate_reg_1[2098])); 
mux_module mux_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4195]),.i2(intermediate_reg_0[4194]),.o(intermediate_reg_1[2097]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4193]),.i2(intermediate_reg_0[4192]),.o(intermediate_reg_1[2096])); 
fsm fsm_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4191]),.i2(intermediate_reg_0[4190]),.o(intermediate_reg_1[2095])); 
fsm fsm_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4189]),.i2(intermediate_reg_0[4188]),.o(intermediate_reg_1[2094])); 
fsm fsm_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4187]),.i2(intermediate_reg_0[4186]),.o(intermediate_reg_1[2093])); 
mux_module mux_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4185]),.i2(intermediate_reg_0[4184]),.o(intermediate_reg_1[2092]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4183]),.i2(intermediate_reg_0[4182]),.o(intermediate_reg_1[2091])); 
mux_module mux_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4181]),.i2(intermediate_reg_0[4180]),.o(intermediate_reg_1[2090]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4179]),.i2(intermediate_reg_0[4178]),.o(intermediate_reg_1[2089])); 
fsm fsm_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4177]),.i2(intermediate_reg_0[4176]),.o(intermediate_reg_1[2088])); 
fsm fsm_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4175]),.i2(intermediate_reg_0[4174]),.o(intermediate_reg_1[2087])); 
mux_module mux_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4173]),.i2(intermediate_reg_0[4172]),.o(intermediate_reg_1[2086]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4171]),.i2(intermediate_reg_0[4170]),.o(intermediate_reg_1[2085])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4169]),.i2(intermediate_reg_0[4168]),.o(intermediate_reg_1[2084]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4167]),.i2(intermediate_reg_0[4166]),.o(intermediate_reg_1[2083])); 
fsm fsm_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4165]),.i2(intermediate_reg_0[4164]),.o(intermediate_reg_1[2082])); 
mux_module mux_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4163]),.i2(intermediate_reg_0[4162]),.o(intermediate_reg_1[2081]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4161]),.i2(intermediate_reg_0[4160]),.o(intermediate_reg_1[2080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4159]),.i2(intermediate_reg_0[4158]),.o(intermediate_reg_1[2079]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4157]),.i2(intermediate_reg_0[4156]),.o(intermediate_reg_1[2078])); 
fsm fsm_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4155]),.i2(intermediate_reg_0[4154]),.o(intermediate_reg_1[2077])); 
mux_module mux_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4153]),.i2(intermediate_reg_0[4152]),.o(intermediate_reg_1[2076]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4151]),.i2(intermediate_reg_0[4150]),.o(intermediate_reg_1[2075]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4149]),.i2(intermediate_reg_0[4148]),.o(intermediate_reg_1[2074])); 
mux_module mux_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4147]),.i2(intermediate_reg_0[4146]),.o(intermediate_reg_1[2073]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4145]),.i2(intermediate_reg_0[4144]),.o(intermediate_reg_1[2072]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4143]),.i2(intermediate_reg_0[4142]),.o(intermediate_reg_1[2071]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4141]),.i2(intermediate_reg_0[4140]),.o(intermediate_reg_1[2070])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4139]),.i2(intermediate_reg_0[4138]),.o(intermediate_reg_1[2069]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4137]),.i2(intermediate_reg_0[4136]),.o(intermediate_reg_1[2068])); 
mux_module mux_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4135]),.i2(intermediate_reg_0[4134]),.o(intermediate_reg_1[2067]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4133]),.i2(intermediate_reg_0[4132]),.o(intermediate_reg_1[2066]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4131]),.i2(intermediate_reg_0[4130]),.o(intermediate_reg_1[2065]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4129]),.i2(intermediate_reg_0[4128]),.o(intermediate_reg_1[2064]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4127]),.i2(intermediate_reg_0[4126]),.o(intermediate_reg_1[2063]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4125]),.i2(intermediate_reg_0[4124]),.o(intermediate_reg_1[2062]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4123]),.i2(intermediate_reg_0[4122]),.o(intermediate_reg_1[2061])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4121]),.i2(intermediate_reg_0[4120]),.o(intermediate_reg_1[2060]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4119]),.i2(intermediate_reg_0[4118]),.o(intermediate_reg_1[2059])); 
fsm fsm_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4117]),.i2(intermediate_reg_0[4116]),.o(intermediate_reg_1[2058])); 
mux_module mux_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4115]),.i2(intermediate_reg_0[4114]),.o(intermediate_reg_1[2057]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4113]),.i2(intermediate_reg_0[4112]),.o(intermediate_reg_1[2056]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4111]),.i2(intermediate_reg_0[4110]),.o(intermediate_reg_1[2055]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4109]),.i2(intermediate_reg_0[4108]),.o(intermediate_reg_1[2054])); 
mux_module mux_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4107]),.i2(intermediate_reg_0[4106]),.o(intermediate_reg_1[2053]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4105]),.i2(intermediate_reg_0[4104]),.o(intermediate_reg_1[2052])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4103]),.i2(intermediate_reg_0[4102]),.o(intermediate_reg_1[2051]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4101]),.i2(intermediate_reg_0[4100]),.o(intermediate_reg_1[2050])); 
mux_module mux_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4099]),.i2(intermediate_reg_0[4098]),.o(intermediate_reg_1[2049]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4097]),.i2(intermediate_reg_0[4096]),.o(intermediate_reg_1[2048]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4095]),.i2(intermediate_reg_0[4094]),.o(intermediate_reg_1[2047])); 
fsm fsm_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4093]),.i2(intermediate_reg_0[4092]),.o(intermediate_reg_1[2046])); 
mux_module mux_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4091]),.i2(intermediate_reg_0[4090]),.o(intermediate_reg_1[2045]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4089]),.i2(intermediate_reg_0[4088]),.o(intermediate_reg_1[2044]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4087]),.i2(intermediate_reg_0[4086]),.o(intermediate_reg_1[2043]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4085]),.i2(intermediate_reg_0[4084]),.o(intermediate_reg_1[2042]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4083]),.i2(intermediate_reg_0[4082]),.o(intermediate_reg_1[2041])); 
fsm fsm_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4081]),.i2(intermediate_reg_0[4080]),.o(intermediate_reg_1[2040])); 
fsm fsm_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4079]),.i2(intermediate_reg_0[4078]),.o(intermediate_reg_1[2039])); 
fsm fsm_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4077]),.i2(intermediate_reg_0[4076]),.o(intermediate_reg_1[2038])); 
mux_module mux_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4075]),.i2(intermediate_reg_0[4074]),.o(intermediate_reg_1[2037]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4073]),.i2(intermediate_reg_0[4072]),.o(intermediate_reg_1[2036])); 
mux_module mux_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4071]),.i2(intermediate_reg_0[4070]),.o(intermediate_reg_1[2035]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4069]),.i2(intermediate_reg_0[4068]),.o(intermediate_reg_1[2034]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4067]),.i2(intermediate_reg_0[4066]),.o(intermediate_reg_1[2033])); 
fsm fsm_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4065]),.i2(intermediate_reg_0[4064]),.o(intermediate_reg_1[2032])); 
mux_module mux_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4063]),.i2(intermediate_reg_0[4062]),.o(intermediate_reg_1[2031]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4061]),.i2(intermediate_reg_0[4060]),.o(intermediate_reg_1[2030]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4059]),.i2(intermediate_reg_0[4058]),.o(intermediate_reg_1[2029])); 
fsm fsm_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4057]),.i2(intermediate_reg_0[4056]),.o(intermediate_reg_1[2028])); 
mux_module mux_module_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4055]),.i2(intermediate_reg_0[4054]),.o(intermediate_reg_1[2027]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4053]),.i2(intermediate_reg_0[4052]),.o(intermediate_reg_1[2026])); 
mux_module mux_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4051]),.i2(intermediate_reg_0[4050]),.o(intermediate_reg_1[2025]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4049]),.i2(intermediate_reg_0[4048]),.o(intermediate_reg_1[2024])); 
fsm fsm_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4047]),.i2(intermediate_reg_0[4046]),.o(intermediate_reg_1[2023])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4045]),.i2(intermediate_reg_0[4044]),.o(intermediate_reg_1[2022]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4043]),.i2(intermediate_reg_0[4042]),.o(intermediate_reg_1[2021])); 
fsm fsm_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4041]),.i2(intermediate_reg_0[4040]),.o(intermediate_reg_1[2020])); 
mux_module mux_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4039]),.i2(intermediate_reg_0[4038]),.o(intermediate_reg_1[2019]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4037]),.i2(intermediate_reg_0[4036]),.o(intermediate_reg_1[2018])); 
mux_module mux_module_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4035]),.i2(intermediate_reg_0[4034]),.o(intermediate_reg_1[2017]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4033]),.i2(intermediate_reg_0[4032]),.o(intermediate_reg_1[2016]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4031]),.i2(intermediate_reg_0[4030]),.o(intermediate_reg_1[2015])); 
fsm fsm_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4029]),.i2(intermediate_reg_0[4028]),.o(intermediate_reg_1[2014])); 
mux_module mux_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4027]),.i2(intermediate_reg_0[4026]),.o(intermediate_reg_1[2013]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4025]),.i2(intermediate_reg_0[4024]),.o(intermediate_reg_1[2012]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4023]),.i2(intermediate_reg_0[4022]),.o(intermediate_reg_1[2011])); 
mux_module mux_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4021]),.i2(intermediate_reg_0[4020]),.o(intermediate_reg_1[2010]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4019]),.i2(intermediate_reg_0[4018]),.o(intermediate_reg_1[2009])); 
mux_module mux_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4017]),.i2(intermediate_reg_0[4016]),.o(intermediate_reg_1[2008]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4015]),.i2(intermediate_reg_0[4014]),.o(intermediate_reg_1[2007])); 
mux_module mux_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4013]),.i2(intermediate_reg_0[4012]),.o(intermediate_reg_1[2006]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4011]),.i2(intermediate_reg_0[4010]),.o(intermediate_reg_1[2005])); 
fsm fsm_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4009]),.i2(intermediate_reg_0[4008]),.o(intermediate_reg_1[2004])); 
fsm fsm_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4007]),.i2(intermediate_reg_0[4006]),.o(intermediate_reg_1[2003])); 
mux_module mux_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4005]),.i2(intermediate_reg_0[4004]),.o(intermediate_reg_1[2002]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4003]),.i2(intermediate_reg_0[4002]),.o(intermediate_reg_1[2001])); 
mux_module mux_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4001]),.i2(intermediate_reg_0[4000]),.o(intermediate_reg_1[2000]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3999]),.i2(intermediate_reg_0[3998]),.o(intermediate_reg_1[1999]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3997]),.i2(intermediate_reg_0[3996]),.o(intermediate_reg_1[1998])); 
mux_module mux_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3995]),.i2(intermediate_reg_0[3994]),.o(intermediate_reg_1[1997]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3993]),.i2(intermediate_reg_0[3992]),.o(intermediate_reg_1[1996])); 
fsm fsm_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3991]),.i2(intermediate_reg_0[3990]),.o(intermediate_reg_1[1995])); 
mux_module mux_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3989]),.i2(intermediate_reg_0[3988]),.o(intermediate_reg_1[1994]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3987]),.i2(intermediate_reg_0[3986]),.o(intermediate_reg_1[1993]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3985]),.i2(intermediate_reg_0[3984]),.o(intermediate_reg_1[1992])); 
mux_module mux_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3983]),.i2(intermediate_reg_0[3982]),.o(intermediate_reg_1[1991]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3981]),.i2(intermediate_reg_0[3980]),.o(intermediate_reg_1[1990])); 
fsm fsm_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3979]),.i2(intermediate_reg_0[3978]),.o(intermediate_reg_1[1989])); 
mux_module mux_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3977]),.i2(intermediate_reg_0[3976]),.o(intermediate_reg_1[1988]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3975]),.i2(intermediate_reg_0[3974]),.o(intermediate_reg_1[1987]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3973]),.i2(intermediate_reg_0[3972]),.o(intermediate_reg_1[1986]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3971]),.i2(intermediate_reg_0[3970]),.o(intermediate_reg_1[1985])); 
fsm fsm_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3969]),.i2(intermediate_reg_0[3968]),.o(intermediate_reg_1[1984])); 
fsm fsm_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3967]),.i2(intermediate_reg_0[3966]),.o(intermediate_reg_1[1983])); 
mux_module mux_module_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3965]),.i2(intermediate_reg_0[3964]),.o(intermediate_reg_1[1982]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3963]),.i2(intermediate_reg_0[3962]),.o(intermediate_reg_1[1981])); 
fsm fsm_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3961]),.i2(intermediate_reg_0[3960]),.o(intermediate_reg_1[1980])); 
fsm fsm_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3959]),.i2(intermediate_reg_0[3958]),.o(intermediate_reg_1[1979])); 
mux_module mux_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3957]),.i2(intermediate_reg_0[3956]),.o(intermediate_reg_1[1978]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3955]),.i2(intermediate_reg_0[3954]),.o(intermediate_reg_1[1977])); 
mux_module mux_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3953]),.i2(intermediate_reg_0[3952]),.o(intermediate_reg_1[1976]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3951]),.i2(intermediate_reg_0[3950]),.o(intermediate_reg_1[1975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3949]),.i2(intermediate_reg_0[3948]),.o(intermediate_reg_1[1974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3947]),.i2(intermediate_reg_0[3946]),.o(intermediate_reg_1[1973]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3945]),.i2(intermediate_reg_0[3944]),.o(intermediate_reg_1[1972]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3943]),.i2(intermediate_reg_0[3942]),.o(intermediate_reg_1[1971]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3941]),.i2(intermediate_reg_0[3940]),.o(intermediate_reg_1[1970])); 
fsm fsm_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3939]),.i2(intermediate_reg_0[3938]),.o(intermediate_reg_1[1969])); 
fsm fsm_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3937]),.i2(intermediate_reg_0[3936]),.o(intermediate_reg_1[1968])); 
fsm fsm_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3935]),.i2(intermediate_reg_0[3934]),.o(intermediate_reg_1[1967])); 
fsm fsm_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3933]),.i2(intermediate_reg_0[3932]),.o(intermediate_reg_1[1966])); 
fsm fsm_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3931]),.i2(intermediate_reg_0[3930]),.o(intermediate_reg_1[1965])); 
fsm fsm_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3929]),.i2(intermediate_reg_0[3928]),.o(intermediate_reg_1[1964])); 
mux_module mux_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3927]),.i2(intermediate_reg_0[3926]),.o(intermediate_reg_1[1963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3925]),.i2(intermediate_reg_0[3924]),.o(intermediate_reg_1[1962]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3923]),.i2(intermediate_reg_0[3922]),.o(intermediate_reg_1[1961]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3921]),.i2(intermediate_reg_0[3920]),.o(intermediate_reg_1[1960]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3919]),.i2(intermediate_reg_0[3918]),.o(intermediate_reg_1[1959])); 
mux_module mux_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3917]),.i2(intermediate_reg_0[3916]),.o(intermediate_reg_1[1958]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3915]),.i2(intermediate_reg_0[3914]),.o(intermediate_reg_1[1957]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3913]),.i2(intermediate_reg_0[3912]),.o(intermediate_reg_1[1956])); 
mux_module mux_module_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3911]),.i2(intermediate_reg_0[3910]),.o(intermediate_reg_1[1955]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3909]),.i2(intermediate_reg_0[3908]),.o(intermediate_reg_1[1954]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3907]),.i2(intermediate_reg_0[3906]),.o(intermediate_reg_1[1953]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3905]),.i2(intermediate_reg_0[3904]),.o(intermediate_reg_1[1952]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3903]),.i2(intermediate_reg_0[3902]),.o(intermediate_reg_1[1951]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3901]),.i2(intermediate_reg_0[3900]),.o(intermediate_reg_1[1950])); 
mux_module mux_module_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3899]),.i2(intermediate_reg_0[3898]),.o(intermediate_reg_1[1949]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3897]),.i2(intermediate_reg_0[3896]),.o(intermediate_reg_1[1948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3895]),.i2(intermediate_reg_0[3894]),.o(intermediate_reg_1[1947]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3893]),.i2(intermediate_reg_0[3892]),.o(intermediate_reg_1[1946])); 
fsm fsm_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3891]),.i2(intermediate_reg_0[3890]),.o(intermediate_reg_1[1945])); 
fsm fsm_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3889]),.i2(intermediate_reg_0[3888]),.o(intermediate_reg_1[1944])); 
fsm fsm_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3887]),.i2(intermediate_reg_0[3886]),.o(intermediate_reg_1[1943])); 
fsm fsm_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3885]),.i2(intermediate_reg_0[3884]),.o(intermediate_reg_1[1942])); 
fsm fsm_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3883]),.i2(intermediate_reg_0[3882]),.o(intermediate_reg_1[1941])); 
mux_module mux_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3881]),.i2(intermediate_reg_0[3880]),.o(intermediate_reg_1[1940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3879]),.i2(intermediate_reg_0[3878]),.o(intermediate_reg_1[1939]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3877]),.i2(intermediate_reg_0[3876]),.o(intermediate_reg_1[1938])); 
fsm fsm_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3875]),.i2(intermediate_reg_0[3874]),.o(intermediate_reg_1[1937])); 
mux_module mux_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3873]),.i2(intermediate_reg_0[3872]),.o(intermediate_reg_1[1936]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3871]),.i2(intermediate_reg_0[3870]),.o(intermediate_reg_1[1935])); 
fsm fsm_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3869]),.i2(intermediate_reg_0[3868]),.o(intermediate_reg_1[1934])); 
fsm fsm_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3867]),.i2(intermediate_reg_0[3866]),.o(intermediate_reg_1[1933])); 
mux_module mux_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3865]),.i2(intermediate_reg_0[3864]),.o(intermediate_reg_1[1932]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3863]),.i2(intermediate_reg_0[3862]),.o(intermediate_reg_1[1931])); 
mux_module mux_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3861]),.i2(intermediate_reg_0[3860]),.o(intermediate_reg_1[1930]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3859]),.i2(intermediate_reg_0[3858]),.o(intermediate_reg_1[1929])); 
mux_module mux_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3857]),.i2(intermediate_reg_0[3856]),.o(intermediate_reg_1[1928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3855]),.i2(intermediate_reg_0[3854]),.o(intermediate_reg_1[1927]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3853]),.i2(intermediate_reg_0[3852]),.o(intermediate_reg_1[1926]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3851]),.i2(intermediate_reg_0[3850]),.o(intermediate_reg_1[1925])); 
fsm fsm_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3849]),.i2(intermediate_reg_0[3848]),.o(intermediate_reg_1[1924])); 
fsm fsm_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3847]),.i2(intermediate_reg_0[3846]),.o(intermediate_reg_1[1923])); 
fsm fsm_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3845]),.i2(intermediate_reg_0[3844]),.o(intermediate_reg_1[1922])); 
mux_module mux_module_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3843]),.i2(intermediate_reg_0[3842]),.o(intermediate_reg_1[1921]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3841]),.i2(intermediate_reg_0[3840]),.o(intermediate_reg_1[1920])); 
fsm fsm_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3839]),.i2(intermediate_reg_0[3838]),.o(intermediate_reg_1[1919])); 
mux_module mux_module_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3837]),.i2(intermediate_reg_0[3836]),.o(intermediate_reg_1[1918]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3835]),.i2(intermediate_reg_0[3834]),.o(intermediate_reg_1[1917])); 
fsm fsm_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3833]),.i2(intermediate_reg_0[3832]),.o(intermediate_reg_1[1916])); 
mux_module mux_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3831]),.i2(intermediate_reg_0[3830]),.o(intermediate_reg_1[1915]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3829]),.i2(intermediate_reg_0[3828]),.o(intermediate_reg_1[1914])); 
mux_module mux_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3827]),.i2(intermediate_reg_0[3826]),.o(intermediate_reg_1[1913]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3825]),.i2(intermediate_reg_0[3824]),.o(intermediate_reg_1[1912])); 
fsm fsm_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3823]),.i2(intermediate_reg_0[3822]),.o(intermediate_reg_1[1911])); 
fsm fsm_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3821]),.i2(intermediate_reg_0[3820]),.o(intermediate_reg_1[1910])); 
mux_module mux_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3819]),.i2(intermediate_reg_0[3818]),.o(intermediate_reg_1[1909]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3817]),.i2(intermediate_reg_0[3816]),.o(intermediate_reg_1[1908]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3815]),.i2(intermediate_reg_0[3814]),.o(intermediate_reg_1[1907]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3813]),.i2(intermediate_reg_0[3812]),.o(intermediate_reg_1[1906])); 
mux_module mux_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3811]),.i2(intermediate_reg_0[3810]),.o(intermediate_reg_1[1905]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3809]),.i2(intermediate_reg_0[3808]),.o(intermediate_reg_1[1904])); 
fsm fsm_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3807]),.i2(intermediate_reg_0[3806]),.o(intermediate_reg_1[1903])); 
fsm fsm_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3805]),.i2(intermediate_reg_0[3804]),.o(intermediate_reg_1[1902])); 
fsm fsm_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3803]),.i2(intermediate_reg_0[3802]),.o(intermediate_reg_1[1901])); 
mux_module mux_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3801]),.i2(intermediate_reg_0[3800]),.o(intermediate_reg_1[1900]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3799]),.i2(intermediate_reg_0[3798]),.o(intermediate_reg_1[1899]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3797]),.i2(intermediate_reg_0[3796]),.o(intermediate_reg_1[1898]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3795]),.i2(intermediate_reg_0[3794]),.o(intermediate_reg_1[1897])); 
fsm fsm_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3793]),.i2(intermediate_reg_0[3792]),.o(intermediate_reg_1[1896])); 
fsm fsm_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3791]),.i2(intermediate_reg_0[3790]),.o(intermediate_reg_1[1895])); 
mux_module mux_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3789]),.i2(intermediate_reg_0[3788]),.o(intermediate_reg_1[1894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3787]),.i2(intermediate_reg_0[3786]),.o(intermediate_reg_1[1893]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3785]),.i2(intermediate_reg_0[3784]),.o(intermediate_reg_1[1892])); 
mux_module mux_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3783]),.i2(intermediate_reg_0[3782]),.o(intermediate_reg_1[1891]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3781]),.i2(intermediate_reg_0[3780]),.o(intermediate_reg_1[1890]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3779]),.i2(intermediate_reg_0[3778]),.o(intermediate_reg_1[1889])); 
mux_module mux_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3777]),.i2(intermediate_reg_0[3776]),.o(intermediate_reg_1[1888]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3775]),.i2(intermediate_reg_0[3774]),.o(intermediate_reg_1[1887])); 
mux_module mux_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3773]),.i2(intermediate_reg_0[3772]),.o(intermediate_reg_1[1886]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3771]),.i2(intermediate_reg_0[3770]),.o(intermediate_reg_1[1885])); 
fsm fsm_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3769]),.i2(intermediate_reg_0[3768]),.o(intermediate_reg_1[1884])); 
mux_module mux_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3767]),.i2(intermediate_reg_0[3766]),.o(intermediate_reg_1[1883]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3765]),.i2(intermediate_reg_0[3764]),.o(intermediate_reg_1[1882]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3763]),.i2(intermediate_reg_0[3762]),.o(intermediate_reg_1[1881]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3761]),.i2(intermediate_reg_0[3760]),.o(intermediate_reg_1[1880])); 
mux_module mux_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3759]),.i2(intermediate_reg_0[3758]),.o(intermediate_reg_1[1879]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3757]),.i2(intermediate_reg_0[3756]),.o(intermediate_reg_1[1878])); 
fsm fsm_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3755]),.i2(intermediate_reg_0[3754]),.o(intermediate_reg_1[1877])); 
fsm fsm_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3753]),.i2(intermediate_reg_0[3752]),.o(intermediate_reg_1[1876])); 
mux_module mux_module_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3751]),.i2(intermediate_reg_0[3750]),.o(intermediate_reg_1[1875]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3749]),.i2(intermediate_reg_0[3748]),.o(intermediate_reg_1[1874]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3747]),.i2(intermediate_reg_0[3746]),.o(intermediate_reg_1[1873])); 
fsm fsm_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3745]),.i2(intermediate_reg_0[3744]),.o(intermediate_reg_1[1872])); 
mux_module mux_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3743]),.i2(intermediate_reg_0[3742]),.o(intermediate_reg_1[1871]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3741]),.i2(intermediate_reg_0[3740]),.o(intermediate_reg_1[1870])); 
fsm fsm_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3739]),.i2(intermediate_reg_0[3738]),.o(intermediate_reg_1[1869])); 
fsm fsm_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3737]),.i2(intermediate_reg_0[3736]),.o(intermediate_reg_1[1868])); 
fsm fsm_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3735]),.i2(intermediate_reg_0[3734]),.o(intermediate_reg_1[1867])); 
mux_module mux_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3733]),.i2(intermediate_reg_0[3732]),.o(intermediate_reg_1[1866]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3731]),.i2(intermediate_reg_0[3730]),.o(intermediate_reg_1[1865])); 
fsm fsm_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3729]),.i2(intermediate_reg_0[3728]),.o(intermediate_reg_1[1864])); 
mux_module mux_module_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3727]),.i2(intermediate_reg_0[3726]),.o(intermediate_reg_1[1863]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3725]),.i2(intermediate_reg_0[3724]),.o(intermediate_reg_1[1862])); 
mux_module mux_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3723]),.i2(intermediate_reg_0[3722]),.o(intermediate_reg_1[1861]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3721]),.i2(intermediate_reg_0[3720]),.o(intermediate_reg_1[1860]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3719]),.i2(intermediate_reg_0[3718]),.o(intermediate_reg_1[1859])); 
fsm fsm_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3717]),.i2(intermediate_reg_0[3716]),.o(intermediate_reg_1[1858])); 
mux_module mux_module_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3715]),.i2(intermediate_reg_0[3714]),.o(intermediate_reg_1[1857]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3713]),.i2(intermediate_reg_0[3712]),.o(intermediate_reg_1[1856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3711]),.i2(intermediate_reg_0[3710]),.o(intermediate_reg_1[1855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3709]),.i2(intermediate_reg_0[3708]),.o(intermediate_reg_1[1854]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3707]),.i2(intermediate_reg_0[3706]),.o(intermediate_reg_1[1853]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3705]),.i2(intermediate_reg_0[3704]),.o(intermediate_reg_1[1852]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3703]),.i2(intermediate_reg_0[3702]),.o(intermediate_reg_1[1851])); 
fsm fsm_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3701]),.i2(intermediate_reg_0[3700]),.o(intermediate_reg_1[1850])); 
mux_module mux_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3699]),.i2(intermediate_reg_0[3698]),.o(intermediate_reg_1[1849]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3697]),.i2(intermediate_reg_0[3696]),.o(intermediate_reg_1[1848])); 
fsm fsm_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3695]),.i2(intermediate_reg_0[3694]),.o(intermediate_reg_1[1847])); 
fsm fsm_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3693]),.i2(intermediate_reg_0[3692]),.o(intermediate_reg_1[1846])); 
mux_module mux_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3691]),.i2(intermediate_reg_0[3690]),.o(intermediate_reg_1[1845]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3689]),.i2(intermediate_reg_0[3688]),.o(intermediate_reg_1[1844])); 
mux_module mux_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3687]),.i2(intermediate_reg_0[3686]),.o(intermediate_reg_1[1843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3685]),.i2(intermediate_reg_0[3684]),.o(intermediate_reg_1[1842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3683]),.i2(intermediate_reg_0[3682]),.o(intermediate_reg_1[1841]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3681]),.i2(intermediate_reg_0[3680]),.o(intermediate_reg_1[1840])); 
mux_module mux_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3679]),.i2(intermediate_reg_0[3678]),.o(intermediate_reg_1[1839]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3677]),.i2(intermediate_reg_0[3676]),.o(intermediate_reg_1[1838])); 
fsm fsm_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3675]),.i2(intermediate_reg_0[3674]),.o(intermediate_reg_1[1837])); 
fsm fsm_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3673]),.i2(intermediate_reg_0[3672]),.o(intermediate_reg_1[1836])); 
fsm fsm_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3671]),.i2(intermediate_reg_0[3670]),.o(intermediate_reg_1[1835])); 
mux_module mux_module_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3669]),.i2(intermediate_reg_0[3668]),.o(intermediate_reg_1[1834]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3667]),.i2(intermediate_reg_0[3666]),.o(intermediate_reg_1[1833])); 
fsm fsm_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3665]),.i2(intermediate_reg_0[3664]),.o(intermediate_reg_1[1832])); 
mux_module mux_module_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3663]),.i2(intermediate_reg_0[3662]),.o(intermediate_reg_1[1831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3661]),.i2(intermediate_reg_0[3660]),.o(intermediate_reg_1[1830]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3659]),.i2(intermediate_reg_0[3658]),.o(intermediate_reg_1[1829])); 
fsm fsm_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3657]),.i2(intermediate_reg_0[3656]),.o(intermediate_reg_1[1828])); 
fsm fsm_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3655]),.i2(intermediate_reg_0[3654]),.o(intermediate_reg_1[1827])); 
fsm fsm_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3653]),.i2(intermediate_reg_0[3652]),.o(intermediate_reg_1[1826])); 
mux_module mux_module_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3651]),.i2(intermediate_reg_0[3650]),.o(intermediate_reg_1[1825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3649]),.i2(intermediate_reg_0[3648]),.o(intermediate_reg_1[1824]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3647]),.i2(intermediate_reg_0[3646]),.o(intermediate_reg_1[1823])); 
fsm fsm_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3645]),.i2(intermediate_reg_0[3644]),.o(intermediate_reg_1[1822])); 
mux_module mux_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3643]),.i2(intermediate_reg_0[3642]),.o(intermediate_reg_1[1821]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3641]),.i2(intermediate_reg_0[3640]),.o(intermediate_reg_1[1820])); 
mux_module mux_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3639]),.i2(intermediate_reg_0[3638]),.o(intermediate_reg_1[1819]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3637]),.i2(intermediate_reg_0[3636]),.o(intermediate_reg_1[1818]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3635]),.i2(intermediate_reg_0[3634]),.o(intermediate_reg_1[1817])); 
mux_module mux_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3633]),.i2(intermediate_reg_0[3632]),.o(intermediate_reg_1[1816]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3631]),.i2(intermediate_reg_0[3630]),.o(intermediate_reg_1[1815])); 
mux_module mux_module_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3629]),.i2(intermediate_reg_0[3628]),.o(intermediate_reg_1[1814]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3627]),.i2(intermediate_reg_0[3626]),.o(intermediate_reg_1[1813])); 
mux_module mux_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3625]),.i2(intermediate_reg_0[3624]),.o(intermediate_reg_1[1812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3623]),.i2(intermediate_reg_0[3622]),.o(intermediate_reg_1[1811]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3621]),.i2(intermediate_reg_0[3620]),.o(intermediate_reg_1[1810])); 
fsm fsm_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3619]),.i2(intermediate_reg_0[3618]),.o(intermediate_reg_1[1809])); 
mux_module mux_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3617]),.i2(intermediate_reg_0[3616]),.o(intermediate_reg_1[1808]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3615]),.i2(intermediate_reg_0[3614]),.o(intermediate_reg_1[1807])); 
fsm fsm_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3613]),.i2(intermediate_reg_0[3612]),.o(intermediate_reg_1[1806])); 
mux_module mux_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3611]),.i2(intermediate_reg_0[3610]),.o(intermediate_reg_1[1805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3609]),.i2(intermediate_reg_0[3608]),.o(intermediate_reg_1[1804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3607]),.i2(intermediate_reg_0[3606]),.o(intermediate_reg_1[1803]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3605]),.i2(intermediate_reg_0[3604]),.o(intermediate_reg_1[1802]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3603]),.i2(intermediate_reg_0[3602]),.o(intermediate_reg_1[1801])); 
fsm fsm_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3601]),.i2(intermediate_reg_0[3600]),.o(intermediate_reg_1[1800])); 
mux_module mux_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3599]),.i2(intermediate_reg_0[3598]),.o(intermediate_reg_1[1799]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3597]),.i2(intermediate_reg_0[3596]),.o(intermediate_reg_1[1798]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3595]),.i2(intermediate_reg_0[3594]),.o(intermediate_reg_1[1797]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3593]),.i2(intermediate_reg_0[3592]),.o(intermediate_reg_1[1796]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3591]),.i2(intermediate_reg_0[3590]),.o(intermediate_reg_1[1795])); 
fsm fsm_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3589]),.i2(intermediate_reg_0[3588]),.o(intermediate_reg_1[1794])); 
mux_module mux_module_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3587]),.i2(intermediate_reg_0[3586]),.o(intermediate_reg_1[1793]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3585]),.i2(intermediate_reg_0[3584]),.o(intermediate_reg_1[1792]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3583]),.i2(intermediate_reg_0[3582]),.o(intermediate_reg_1[1791]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3581]),.i2(intermediate_reg_0[3580]),.o(intermediate_reg_1[1790])); 
fsm fsm_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3579]),.i2(intermediate_reg_0[3578]),.o(intermediate_reg_1[1789])); 
fsm fsm_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3577]),.i2(intermediate_reg_0[3576]),.o(intermediate_reg_1[1788])); 
fsm fsm_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3575]),.i2(intermediate_reg_0[3574]),.o(intermediate_reg_1[1787])); 
mux_module mux_module_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3573]),.i2(intermediate_reg_0[3572]),.o(intermediate_reg_1[1786]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3571]),.i2(intermediate_reg_0[3570]),.o(intermediate_reg_1[1785]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3569]),.i2(intermediate_reg_0[3568]),.o(intermediate_reg_1[1784])); 
mux_module mux_module_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3567]),.i2(intermediate_reg_0[3566]),.o(intermediate_reg_1[1783]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3565]),.i2(intermediate_reg_0[3564]),.o(intermediate_reg_1[1782]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3563]),.i2(intermediate_reg_0[3562]),.o(intermediate_reg_1[1781])); 
fsm fsm_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3561]),.i2(intermediate_reg_0[3560]),.o(intermediate_reg_1[1780])); 
mux_module mux_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3559]),.i2(intermediate_reg_0[3558]),.o(intermediate_reg_1[1779]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3557]),.i2(intermediate_reg_0[3556]),.o(intermediate_reg_1[1778]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3555]),.i2(intermediate_reg_0[3554]),.o(intermediate_reg_1[1777]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3553]),.i2(intermediate_reg_0[3552]),.o(intermediate_reg_1[1776])); 
mux_module mux_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3551]),.i2(intermediate_reg_0[3550]),.o(intermediate_reg_1[1775]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3549]),.i2(intermediate_reg_0[3548]),.o(intermediate_reg_1[1774])); 
mux_module mux_module_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3547]),.i2(intermediate_reg_0[3546]),.o(intermediate_reg_1[1773]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3545]),.i2(intermediate_reg_0[3544]),.o(intermediate_reg_1[1772]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3543]),.i2(intermediate_reg_0[3542]),.o(intermediate_reg_1[1771])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3541]),.i2(intermediate_reg_0[3540]),.o(intermediate_reg_1[1770]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3539]),.i2(intermediate_reg_0[3538]),.o(intermediate_reg_1[1769])); 
mux_module mux_module_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3537]),.i2(intermediate_reg_0[3536]),.o(intermediate_reg_1[1768]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3535]),.i2(intermediate_reg_0[3534]),.o(intermediate_reg_1[1767]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3533]),.i2(intermediate_reg_0[3532]),.o(intermediate_reg_1[1766]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3531]),.i2(intermediate_reg_0[3530]),.o(intermediate_reg_1[1765])); 
mux_module mux_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3529]),.i2(intermediate_reg_0[3528]),.o(intermediate_reg_1[1764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3527]),.i2(intermediate_reg_0[3526]),.o(intermediate_reg_1[1763]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3525]),.i2(intermediate_reg_0[3524]),.o(intermediate_reg_1[1762])); 
mux_module mux_module_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3523]),.i2(intermediate_reg_0[3522]),.o(intermediate_reg_1[1761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3521]),.i2(intermediate_reg_0[3520]),.o(intermediate_reg_1[1760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3519]),.i2(intermediate_reg_0[3518]),.o(intermediate_reg_1[1759]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3517]),.i2(intermediate_reg_0[3516]),.o(intermediate_reg_1[1758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3515]),.i2(intermediate_reg_0[3514]),.o(intermediate_reg_1[1757]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3513]),.i2(intermediate_reg_0[3512]),.o(intermediate_reg_1[1756]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3511]),.i2(intermediate_reg_0[3510]),.o(intermediate_reg_1[1755])); 
mux_module mux_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3509]),.i2(intermediate_reg_0[3508]),.o(intermediate_reg_1[1754]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3507]),.i2(intermediate_reg_0[3506]),.o(intermediate_reg_1[1753])); 
fsm fsm_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3505]),.i2(intermediate_reg_0[3504]),.o(intermediate_reg_1[1752])); 
mux_module mux_module_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3503]),.i2(intermediate_reg_0[3502]),.o(intermediate_reg_1[1751]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3501]),.i2(intermediate_reg_0[3500]),.o(intermediate_reg_1[1750]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3499]),.i2(intermediate_reg_0[3498]),.o(intermediate_reg_1[1749])); 
fsm fsm_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3497]),.i2(intermediate_reg_0[3496]),.o(intermediate_reg_1[1748])); 
mux_module mux_module_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3495]),.i2(intermediate_reg_0[3494]),.o(intermediate_reg_1[1747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3493]),.i2(intermediate_reg_0[3492]),.o(intermediate_reg_1[1746]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3491]),.i2(intermediate_reg_0[3490]),.o(intermediate_reg_1[1745])); 
fsm fsm_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3489]),.i2(intermediate_reg_0[3488]),.o(intermediate_reg_1[1744])); 
mux_module mux_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3487]),.i2(intermediate_reg_0[3486]),.o(intermediate_reg_1[1743]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3485]),.i2(intermediate_reg_0[3484]),.o(intermediate_reg_1[1742])); 
fsm fsm_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3483]),.i2(intermediate_reg_0[3482]),.o(intermediate_reg_1[1741])); 
fsm fsm_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3481]),.i2(intermediate_reg_0[3480]),.o(intermediate_reg_1[1740])); 
fsm fsm_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3479]),.i2(intermediate_reg_0[3478]),.o(intermediate_reg_1[1739])); 
fsm fsm_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3477]),.i2(intermediate_reg_0[3476]),.o(intermediate_reg_1[1738])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3475]),.i2(intermediate_reg_0[3474]),.o(intermediate_reg_1[1737]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3473]),.i2(intermediate_reg_0[3472]),.o(intermediate_reg_1[1736])); 
fsm fsm_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3471]),.i2(intermediate_reg_0[3470]),.o(intermediate_reg_1[1735])); 
fsm fsm_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3469]),.i2(intermediate_reg_0[3468]),.o(intermediate_reg_1[1734])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3467]),.i2(intermediate_reg_0[3466]),.o(intermediate_reg_1[1733]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3465]),.i2(intermediate_reg_0[3464]),.o(intermediate_reg_1[1732]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3463]),.i2(intermediate_reg_0[3462]),.o(intermediate_reg_1[1731])); 
fsm fsm_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3461]),.i2(intermediate_reg_0[3460]),.o(intermediate_reg_1[1730])); 
mux_module mux_module_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3459]),.i2(intermediate_reg_0[3458]),.o(intermediate_reg_1[1729]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3457]),.i2(intermediate_reg_0[3456]),.o(intermediate_reg_1[1728])); 
mux_module mux_module_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3455]),.i2(intermediate_reg_0[3454]),.o(intermediate_reg_1[1727]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3453]),.i2(intermediate_reg_0[3452]),.o(intermediate_reg_1[1726]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3451]),.i2(intermediate_reg_0[3450]),.o(intermediate_reg_1[1725])); 
mux_module mux_module_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3449]),.i2(intermediate_reg_0[3448]),.o(intermediate_reg_1[1724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3447]),.i2(intermediate_reg_0[3446]),.o(intermediate_reg_1[1723]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3445]),.i2(intermediate_reg_0[3444]),.o(intermediate_reg_1[1722])); 
fsm fsm_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3443]),.i2(intermediate_reg_0[3442]),.o(intermediate_reg_1[1721])); 
fsm fsm_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3441]),.i2(intermediate_reg_0[3440]),.o(intermediate_reg_1[1720])); 
fsm fsm_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3439]),.i2(intermediate_reg_0[3438]),.o(intermediate_reg_1[1719])); 
mux_module mux_module_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3437]),.i2(intermediate_reg_0[3436]),.o(intermediate_reg_1[1718]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3435]),.i2(intermediate_reg_0[3434]),.o(intermediate_reg_1[1717])); 
mux_module mux_module_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3433]),.i2(intermediate_reg_0[3432]),.o(intermediate_reg_1[1716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3431]),.i2(intermediate_reg_0[3430]),.o(intermediate_reg_1[1715]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3429]),.i2(intermediate_reg_0[3428]),.o(intermediate_reg_1[1714])); 
fsm fsm_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3427]),.i2(intermediate_reg_0[3426]),.o(intermediate_reg_1[1713])); 
fsm fsm_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3425]),.i2(intermediate_reg_0[3424]),.o(intermediate_reg_1[1712])); 
mux_module mux_module_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3423]),.i2(intermediate_reg_0[3422]),.o(intermediate_reg_1[1711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3421]),.i2(intermediate_reg_0[3420]),.o(intermediate_reg_1[1710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3419]),.i2(intermediate_reg_0[3418]),.o(intermediate_reg_1[1709]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3417]),.i2(intermediate_reg_0[3416]),.o(intermediate_reg_1[1708]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3415]),.i2(intermediate_reg_0[3414]),.o(intermediate_reg_1[1707])); 
mux_module mux_module_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3413]),.i2(intermediate_reg_0[3412]),.o(intermediate_reg_1[1706]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3411]),.i2(intermediate_reg_0[3410]),.o(intermediate_reg_1[1705]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3409]),.i2(intermediate_reg_0[3408]),.o(intermediate_reg_1[1704])); 
mux_module mux_module_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3407]),.i2(intermediate_reg_0[3406]),.o(intermediate_reg_1[1703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3405]),.i2(intermediate_reg_0[3404]),.o(intermediate_reg_1[1702]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3403]),.i2(intermediate_reg_0[3402]),.o(intermediate_reg_1[1701])); 
mux_module mux_module_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3401]),.i2(intermediate_reg_0[3400]),.o(intermediate_reg_1[1700]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3399]),.i2(intermediate_reg_0[3398]),.o(intermediate_reg_1[1699]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3397]),.i2(intermediate_reg_0[3396]),.o(intermediate_reg_1[1698])); 
mux_module mux_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3395]),.i2(intermediate_reg_0[3394]),.o(intermediate_reg_1[1697]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3393]),.i2(intermediate_reg_0[3392]),.o(intermediate_reg_1[1696])); 
mux_module mux_module_inst_1_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3391]),.i2(intermediate_reg_0[3390]),.o(intermediate_reg_1[1695]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3389]),.i2(intermediate_reg_0[3388]),.o(intermediate_reg_1[1694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3387]),.i2(intermediate_reg_0[3386]),.o(intermediate_reg_1[1693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3385]),.i2(intermediate_reg_0[3384]),.o(intermediate_reg_1[1692]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3383]),.i2(intermediate_reg_0[3382]),.o(intermediate_reg_1[1691])); 
fsm fsm_inst_1_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3381]),.i2(intermediate_reg_0[3380]),.o(intermediate_reg_1[1690])); 
fsm fsm_inst_1_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3379]),.i2(intermediate_reg_0[3378]),.o(intermediate_reg_1[1689])); 
mux_module mux_module_inst_1_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3377]),.i2(intermediate_reg_0[3376]),.o(intermediate_reg_1[1688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3375]),.i2(intermediate_reg_0[3374]),.o(intermediate_reg_1[1687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3373]),.i2(intermediate_reg_0[3372]),.o(intermediate_reg_1[1686]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3371]),.i2(intermediate_reg_0[3370]),.o(intermediate_reg_1[1685])); 
mux_module mux_module_inst_1_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3369]),.i2(intermediate_reg_0[3368]),.o(intermediate_reg_1[1684]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3367]),.i2(intermediate_reg_0[3366]),.o(intermediate_reg_1[1683])); 
fsm fsm_inst_1_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3365]),.i2(intermediate_reg_0[3364]),.o(intermediate_reg_1[1682])); 
fsm fsm_inst_1_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3363]),.i2(intermediate_reg_0[3362]),.o(intermediate_reg_1[1681])); 
fsm fsm_inst_1_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3361]),.i2(intermediate_reg_0[3360]),.o(intermediate_reg_1[1680])); 
mux_module mux_module_inst_1_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3359]),.i2(intermediate_reg_0[3358]),.o(intermediate_reg_1[1679]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3357]),.i2(intermediate_reg_0[3356]),.o(intermediate_reg_1[1678]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3355]),.i2(intermediate_reg_0[3354]),.o(intermediate_reg_1[1677]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3353]),.i2(intermediate_reg_0[3352]),.o(intermediate_reg_1[1676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3351]),.i2(intermediate_reg_0[3350]),.o(intermediate_reg_1[1675]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3349]),.i2(intermediate_reg_0[3348]),.o(intermediate_reg_1[1674])); 
mux_module mux_module_inst_1_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3347]),.i2(intermediate_reg_0[3346]),.o(intermediate_reg_1[1673]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3345]),.i2(intermediate_reg_0[3344]),.o(intermediate_reg_1[1672])); 
mux_module mux_module_inst_1_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3343]),.i2(intermediate_reg_0[3342]),.o(intermediate_reg_1[1671]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3341]),.i2(intermediate_reg_0[3340]),.o(intermediate_reg_1[1670])); 
fsm fsm_inst_1_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3339]),.i2(intermediate_reg_0[3338]),.o(intermediate_reg_1[1669])); 
mux_module mux_module_inst_1_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3337]),.i2(intermediate_reg_0[3336]),.o(intermediate_reg_1[1668]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3335]),.i2(intermediate_reg_0[3334]),.o(intermediate_reg_1[1667])); 
fsm fsm_inst_1_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3333]),.i2(intermediate_reg_0[3332]),.o(intermediate_reg_1[1666])); 
fsm fsm_inst_1_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3331]),.i2(intermediate_reg_0[3330]),.o(intermediate_reg_1[1665])); 
mux_module mux_module_inst_1_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3329]),.i2(intermediate_reg_0[3328]),.o(intermediate_reg_1[1664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3327]),.i2(intermediate_reg_0[3326]),.o(intermediate_reg_1[1663]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3325]),.i2(intermediate_reg_0[3324]),.o(intermediate_reg_1[1662])); 
mux_module mux_module_inst_1_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3323]),.i2(intermediate_reg_0[3322]),.o(intermediate_reg_1[1661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3321]),.i2(intermediate_reg_0[3320]),.o(intermediate_reg_1[1660]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3319]),.i2(intermediate_reg_0[3318]),.o(intermediate_reg_1[1659])); 
fsm fsm_inst_1_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3317]),.i2(intermediate_reg_0[3316]),.o(intermediate_reg_1[1658])); 
fsm fsm_inst_1_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3315]),.i2(intermediate_reg_0[3314]),.o(intermediate_reg_1[1657])); 
fsm fsm_inst_1_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3313]),.i2(intermediate_reg_0[3312]),.o(intermediate_reg_1[1656])); 
fsm fsm_inst_1_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3311]),.i2(intermediate_reg_0[3310]),.o(intermediate_reg_1[1655])); 
fsm fsm_inst_1_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3309]),.i2(intermediate_reg_0[3308]),.o(intermediate_reg_1[1654])); 
fsm fsm_inst_1_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3307]),.i2(intermediate_reg_0[3306]),.o(intermediate_reg_1[1653])); 
mux_module mux_module_inst_1_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3305]),.i2(intermediate_reg_0[3304]),.o(intermediate_reg_1[1652]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3303]),.i2(intermediate_reg_0[3302]),.o(intermediate_reg_1[1651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3301]),.i2(intermediate_reg_0[3300]),.o(intermediate_reg_1[1650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3299]),.i2(intermediate_reg_0[3298]),.o(intermediate_reg_1[1649]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3297]),.i2(intermediate_reg_0[3296]),.o(intermediate_reg_1[1648])); 
fsm fsm_inst_1_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3295]),.i2(intermediate_reg_0[3294]),.o(intermediate_reg_1[1647])); 
mux_module mux_module_inst_1_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3293]),.i2(intermediate_reg_0[3292]),.o(intermediate_reg_1[1646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3291]),.i2(intermediate_reg_0[3290]),.o(intermediate_reg_1[1645]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3289]),.i2(intermediate_reg_0[3288]),.o(intermediate_reg_1[1644]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3287]),.i2(intermediate_reg_0[3286]),.o(intermediate_reg_1[1643])); 
fsm fsm_inst_1_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3285]),.i2(intermediate_reg_0[3284]),.o(intermediate_reg_1[1642])); 
fsm fsm_inst_1_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3283]),.i2(intermediate_reg_0[3282]),.o(intermediate_reg_1[1641])); 
mux_module mux_module_inst_1_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3281]),.i2(intermediate_reg_0[3280]),.o(intermediate_reg_1[1640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3279]),.i2(intermediate_reg_0[3278]),.o(intermediate_reg_1[1639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3277]),.i2(intermediate_reg_0[3276]),.o(intermediate_reg_1[1638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3275]),.i2(intermediate_reg_0[3274]),.o(intermediate_reg_1[1637])); 
mux_module mux_module_inst_1_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3273]),.i2(intermediate_reg_0[3272]),.o(intermediate_reg_1[1636]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3271]),.i2(intermediate_reg_0[3270]),.o(intermediate_reg_1[1635])); 
fsm fsm_inst_1_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3269]),.i2(intermediate_reg_0[3268]),.o(intermediate_reg_1[1634])); 
mux_module mux_module_inst_1_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3267]),.i2(intermediate_reg_0[3266]),.o(intermediate_reg_1[1633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3265]),.i2(intermediate_reg_0[3264]),.o(intermediate_reg_1[1632]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3263]),.i2(intermediate_reg_0[3262]),.o(intermediate_reg_1[1631])); 
fsm fsm_inst_1_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3261]),.i2(intermediate_reg_0[3260]),.o(intermediate_reg_1[1630])); 
fsm fsm_inst_1_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3259]),.i2(intermediate_reg_0[3258]),.o(intermediate_reg_1[1629])); 
mux_module mux_module_inst_1_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3257]),.i2(intermediate_reg_0[3256]),.o(intermediate_reg_1[1628]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3255]),.i2(intermediate_reg_0[3254]),.o(intermediate_reg_1[1627])); 
mux_module mux_module_inst_1_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3253]),.i2(intermediate_reg_0[3252]),.o(intermediate_reg_1[1626]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3251]),.i2(intermediate_reg_0[3250]),.o(intermediate_reg_1[1625]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3249]),.i2(intermediate_reg_0[3248]),.o(intermediate_reg_1[1624]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3247]),.i2(intermediate_reg_0[3246]),.o(intermediate_reg_1[1623])); 
fsm fsm_inst_1_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3245]),.i2(intermediate_reg_0[3244]),.o(intermediate_reg_1[1622])); 
mux_module mux_module_inst_1_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3243]),.i2(intermediate_reg_0[3242]),.o(intermediate_reg_1[1621]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3241]),.i2(intermediate_reg_0[3240]),.o(intermediate_reg_1[1620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3239]),.i2(intermediate_reg_0[3238]),.o(intermediate_reg_1[1619]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3237]),.i2(intermediate_reg_0[3236]),.o(intermediate_reg_1[1618])); 
mux_module mux_module_inst_1_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3235]),.i2(intermediate_reg_0[3234]),.o(intermediate_reg_1[1617]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3233]),.i2(intermediate_reg_0[3232]),.o(intermediate_reg_1[1616])); 
mux_module mux_module_inst_1_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3231]),.i2(intermediate_reg_0[3230]),.o(intermediate_reg_1[1615]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3229]),.i2(intermediate_reg_0[3228]),.o(intermediate_reg_1[1614])); 
fsm fsm_inst_1_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3227]),.i2(intermediate_reg_0[3226]),.o(intermediate_reg_1[1613])); 
fsm fsm_inst_1_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3225]),.i2(intermediate_reg_0[3224]),.o(intermediate_reg_1[1612])); 
fsm fsm_inst_1_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3223]),.i2(intermediate_reg_0[3222]),.o(intermediate_reg_1[1611])); 
fsm fsm_inst_1_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3221]),.i2(intermediate_reg_0[3220]),.o(intermediate_reg_1[1610])); 
fsm fsm_inst_1_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3219]),.i2(intermediate_reg_0[3218]),.o(intermediate_reg_1[1609])); 
fsm fsm_inst_1_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3217]),.i2(intermediate_reg_0[3216]),.o(intermediate_reg_1[1608])); 
fsm fsm_inst_1_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3215]),.i2(intermediate_reg_0[3214]),.o(intermediate_reg_1[1607])); 
fsm fsm_inst_1_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3213]),.i2(intermediate_reg_0[3212]),.o(intermediate_reg_1[1606])); 
mux_module mux_module_inst_1_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3211]),.i2(intermediate_reg_0[3210]),.o(intermediate_reg_1[1605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3209]),.i2(intermediate_reg_0[3208]),.o(intermediate_reg_1[1604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3207]),.i2(intermediate_reg_0[3206]),.o(intermediate_reg_1[1603]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3205]),.i2(intermediate_reg_0[3204]),.o(intermediate_reg_1[1602]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3203]),.i2(intermediate_reg_0[3202]),.o(intermediate_reg_1[1601]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3201]),.i2(intermediate_reg_0[3200]),.o(intermediate_reg_1[1600]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3199]),.i2(intermediate_reg_0[3198]),.o(intermediate_reg_1[1599]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3197]),.i2(intermediate_reg_0[3196]),.o(intermediate_reg_1[1598]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3195]),.i2(intermediate_reg_0[3194]),.o(intermediate_reg_1[1597]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3193]),.i2(intermediate_reg_0[3192]),.o(intermediate_reg_1[1596])); 
mux_module mux_module_inst_1_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3191]),.i2(intermediate_reg_0[3190]),.o(intermediate_reg_1[1595]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3189]),.i2(intermediate_reg_0[3188]),.o(intermediate_reg_1[1594]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3187]),.i2(intermediate_reg_0[3186]),.o(intermediate_reg_1[1593]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3185]),.i2(intermediate_reg_0[3184]),.o(intermediate_reg_1[1592]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3183]),.i2(intermediate_reg_0[3182]),.o(intermediate_reg_1[1591]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3181]),.i2(intermediate_reg_0[3180]),.o(intermediate_reg_1[1590])); 
fsm fsm_inst_1_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3179]),.i2(intermediate_reg_0[3178]),.o(intermediate_reg_1[1589])); 
mux_module mux_module_inst_1_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3177]),.i2(intermediate_reg_0[3176]),.o(intermediate_reg_1[1588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3175]),.i2(intermediate_reg_0[3174]),.o(intermediate_reg_1[1587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3173]),.i2(intermediate_reg_0[3172]),.o(intermediate_reg_1[1586]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3171]),.i2(intermediate_reg_0[3170]),.o(intermediate_reg_1[1585])); 
fsm fsm_inst_1_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3169]),.i2(intermediate_reg_0[3168]),.o(intermediate_reg_1[1584])); 
fsm fsm_inst_1_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3167]),.i2(intermediate_reg_0[3166]),.o(intermediate_reg_1[1583])); 
mux_module mux_module_inst_1_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3165]),.i2(intermediate_reg_0[3164]),.o(intermediate_reg_1[1582]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3163]),.i2(intermediate_reg_0[3162]),.o(intermediate_reg_1[1581]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3161]),.i2(intermediate_reg_0[3160]),.o(intermediate_reg_1[1580]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3159]),.i2(intermediate_reg_0[3158]),.o(intermediate_reg_1[1579]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3157]),.i2(intermediate_reg_0[3156]),.o(intermediate_reg_1[1578])); 
mux_module mux_module_inst_1_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3155]),.i2(intermediate_reg_0[3154]),.o(intermediate_reg_1[1577]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3153]),.i2(intermediate_reg_0[3152]),.o(intermediate_reg_1[1576])); 
fsm fsm_inst_1_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3151]),.i2(intermediate_reg_0[3150]),.o(intermediate_reg_1[1575])); 
fsm fsm_inst_1_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3149]),.i2(intermediate_reg_0[3148]),.o(intermediate_reg_1[1574])); 
fsm fsm_inst_1_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3147]),.i2(intermediate_reg_0[3146]),.o(intermediate_reg_1[1573])); 
fsm fsm_inst_1_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3145]),.i2(intermediate_reg_0[3144]),.o(intermediate_reg_1[1572])); 
fsm fsm_inst_1_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3143]),.i2(intermediate_reg_0[3142]),.o(intermediate_reg_1[1571])); 
fsm fsm_inst_1_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3141]),.i2(intermediate_reg_0[3140]),.o(intermediate_reg_1[1570])); 
fsm fsm_inst_1_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3139]),.i2(intermediate_reg_0[3138]),.o(intermediate_reg_1[1569])); 
mux_module mux_module_inst_1_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3137]),.i2(intermediate_reg_0[3136]),.o(intermediate_reg_1[1568]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3135]),.i2(intermediate_reg_0[3134]),.o(intermediate_reg_1[1567])); 
mux_module mux_module_inst_1_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3133]),.i2(intermediate_reg_0[3132]),.o(intermediate_reg_1[1566]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3131]),.i2(intermediate_reg_0[3130]),.o(intermediate_reg_1[1565])); 
mux_module mux_module_inst_1_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3129]),.i2(intermediate_reg_0[3128]),.o(intermediate_reg_1[1564]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3127]),.i2(intermediate_reg_0[3126]),.o(intermediate_reg_1[1563])); 
fsm fsm_inst_1_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3125]),.i2(intermediate_reg_0[3124]),.o(intermediate_reg_1[1562])); 
fsm fsm_inst_1_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3123]),.i2(intermediate_reg_0[3122]),.o(intermediate_reg_1[1561])); 
mux_module mux_module_inst_1_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3121]),.i2(intermediate_reg_0[3120]),.o(intermediate_reg_1[1560]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3119]),.i2(intermediate_reg_0[3118]),.o(intermediate_reg_1[1559])); 
fsm fsm_inst_1_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3117]),.i2(intermediate_reg_0[3116]),.o(intermediate_reg_1[1558])); 
mux_module mux_module_inst_1_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3115]),.i2(intermediate_reg_0[3114]),.o(intermediate_reg_1[1557]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3113]),.i2(intermediate_reg_0[3112]),.o(intermediate_reg_1[1556]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3111]),.i2(intermediate_reg_0[3110]),.o(intermediate_reg_1[1555])); 
mux_module mux_module_inst_1_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3109]),.i2(intermediate_reg_0[3108]),.o(intermediate_reg_1[1554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3107]),.i2(intermediate_reg_0[3106]),.o(intermediate_reg_1[1553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3105]),.i2(intermediate_reg_0[3104]),.o(intermediate_reg_1[1552]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3103]),.i2(intermediate_reg_0[3102]),.o(intermediate_reg_1[1551])); 
mux_module mux_module_inst_1_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3101]),.i2(intermediate_reg_0[3100]),.o(intermediate_reg_1[1550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3099]),.i2(intermediate_reg_0[3098]),.o(intermediate_reg_1[1549]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3097]),.i2(intermediate_reg_0[3096]),.o(intermediate_reg_1[1548])); 
fsm fsm_inst_1_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3095]),.i2(intermediate_reg_0[3094]),.o(intermediate_reg_1[1547])); 
mux_module mux_module_inst_1_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3093]),.i2(intermediate_reg_0[3092]),.o(intermediate_reg_1[1546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3091]),.i2(intermediate_reg_0[3090]),.o(intermediate_reg_1[1545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3089]),.i2(intermediate_reg_0[3088]),.o(intermediate_reg_1[1544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3087]),.i2(intermediate_reg_0[3086]),.o(intermediate_reg_1[1543]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3085]),.i2(intermediate_reg_0[3084]),.o(intermediate_reg_1[1542]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3083]),.i2(intermediate_reg_0[3082]),.o(intermediate_reg_1[1541])); 
mux_module mux_module_inst_1_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3081]),.i2(intermediate_reg_0[3080]),.o(intermediate_reg_1[1540]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3079]),.i2(intermediate_reg_0[3078]),.o(intermediate_reg_1[1539])); 
mux_module mux_module_inst_1_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3077]),.i2(intermediate_reg_0[3076]),.o(intermediate_reg_1[1538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3075]),.i2(intermediate_reg_0[3074]),.o(intermediate_reg_1[1537]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3073]),.i2(intermediate_reg_0[3072]),.o(intermediate_reg_1[1536])); 
fsm fsm_inst_1_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3071]),.i2(intermediate_reg_0[3070]),.o(intermediate_reg_1[1535])); 
mux_module mux_module_inst_1_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3069]),.i2(intermediate_reg_0[3068]),.o(intermediate_reg_1[1534]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3067]),.i2(intermediate_reg_0[3066]),.o(intermediate_reg_1[1533])); 
fsm fsm_inst_1_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3065]),.i2(intermediate_reg_0[3064]),.o(intermediate_reg_1[1532])); 
fsm fsm_inst_1_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3063]),.i2(intermediate_reg_0[3062]),.o(intermediate_reg_1[1531])); 
mux_module mux_module_inst_1_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3061]),.i2(intermediate_reg_0[3060]),.o(intermediate_reg_1[1530]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3059]),.i2(intermediate_reg_0[3058]),.o(intermediate_reg_1[1529])); 
fsm fsm_inst_1_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3057]),.i2(intermediate_reg_0[3056]),.o(intermediate_reg_1[1528])); 
fsm fsm_inst_1_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3055]),.i2(intermediate_reg_0[3054]),.o(intermediate_reg_1[1527])); 
mux_module mux_module_inst_1_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3053]),.i2(intermediate_reg_0[3052]),.o(intermediate_reg_1[1526]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3051]),.i2(intermediate_reg_0[3050]),.o(intermediate_reg_1[1525])); 
fsm fsm_inst_1_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3049]),.i2(intermediate_reg_0[3048]),.o(intermediate_reg_1[1524])); 
mux_module mux_module_inst_1_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3047]),.i2(intermediate_reg_0[3046]),.o(intermediate_reg_1[1523]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3045]),.i2(intermediate_reg_0[3044]),.o(intermediate_reg_1[1522])); 
mux_module mux_module_inst_1_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3043]),.i2(intermediate_reg_0[3042]),.o(intermediate_reg_1[1521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3041]),.i2(intermediate_reg_0[3040]),.o(intermediate_reg_1[1520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3039]),.i2(intermediate_reg_0[3038]),.o(intermediate_reg_1[1519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3037]),.i2(intermediate_reg_0[3036]),.o(intermediate_reg_1[1518]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3035]),.i2(intermediate_reg_0[3034]),.o(intermediate_reg_1[1517])); 
fsm fsm_inst_1_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3033]),.i2(intermediate_reg_0[3032]),.o(intermediate_reg_1[1516])); 
mux_module mux_module_inst_1_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3031]),.i2(intermediate_reg_0[3030]),.o(intermediate_reg_1[1515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3029]),.i2(intermediate_reg_0[3028]),.o(intermediate_reg_1[1514]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3027]),.i2(intermediate_reg_0[3026]),.o(intermediate_reg_1[1513]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3025]),.i2(intermediate_reg_0[3024]),.o(intermediate_reg_1[1512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3023]),.i2(intermediate_reg_0[3022]),.o(intermediate_reg_1[1511]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3021]),.i2(intermediate_reg_0[3020]),.o(intermediate_reg_1[1510]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3019]),.i2(intermediate_reg_0[3018]),.o(intermediate_reg_1[1509])); 
fsm fsm_inst_1_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3017]),.i2(intermediate_reg_0[3016]),.o(intermediate_reg_1[1508])); 
fsm fsm_inst_1_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3015]),.i2(intermediate_reg_0[3014]),.o(intermediate_reg_1[1507])); 
mux_module mux_module_inst_1_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3013]),.i2(intermediate_reg_0[3012]),.o(intermediate_reg_1[1506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3011]),.i2(intermediate_reg_0[3010]),.o(intermediate_reg_1[1505]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3009]),.i2(intermediate_reg_0[3008]),.o(intermediate_reg_1[1504])); 
mux_module mux_module_inst_1_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3007]),.i2(intermediate_reg_0[3006]),.o(intermediate_reg_1[1503]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3005]),.i2(intermediate_reg_0[3004]),.o(intermediate_reg_1[1502])); 
mux_module mux_module_inst_1_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3003]),.i2(intermediate_reg_0[3002]),.o(intermediate_reg_1[1501]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3001]),.i2(intermediate_reg_0[3000]),.o(intermediate_reg_1[1500]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2999]),.i2(intermediate_reg_0[2998]),.o(intermediate_reg_1[1499])); 
fsm fsm_inst_1_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2997]),.i2(intermediate_reg_0[2996]),.o(intermediate_reg_1[1498])); 
mux_module mux_module_inst_1_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2995]),.i2(intermediate_reg_0[2994]),.o(intermediate_reg_1[1497]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2993]),.i2(intermediate_reg_0[2992]),.o(intermediate_reg_1[1496])); 
fsm fsm_inst_1_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2991]),.i2(intermediate_reg_0[2990]),.o(intermediate_reg_1[1495])); 
mux_module mux_module_inst_1_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2989]),.i2(intermediate_reg_0[2988]),.o(intermediate_reg_1[1494]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2987]),.i2(intermediate_reg_0[2986]),.o(intermediate_reg_1[1493])); 
mux_module mux_module_inst_1_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2985]),.i2(intermediate_reg_0[2984]),.o(intermediate_reg_1[1492]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2983]),.i2(intermediate_reg_0[2982]),.o(intermediate_reg_1[1491]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2981]),.i2(intermediate_reg_0[2980]),.o(intermediate_reg_1[1490]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2979]),.i2(intermediate_reg_0[2978]),.o(intermediate_reg_1[1489]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2977]),.i2(intermediate_reg_0[2976]),.o(intermediate_reg_1[1488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2975]),.i2(intermediate_reg_0[2974]),.o(intermediate_reg_1[1487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2973]),.i2(intermediate_reg_0[2972]),.o(intermediate_reg_1[1486]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2971]),.i2(intermediate_reg_0[2970]),.o(intermediate_reg_1[1485])); 
mux_module mux_module_inst_1_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2969]),.i2(intermediate_reg_0[2968]),.o(intermediate_reg_1[1484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2967]),.i2(intermediate_reg_0[2966]),.o(intermediate_reg_1[1483]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2965]),.i2(intermediate_reg_0[2964]),.o(intermediate_reg_1[1482]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2963]),.i2(intermediate_reg_0[2962]),.o(intermediate_reg_1[1481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2961]),.i2(intermediate_reg_0[2960]),.o(intermediate_reg_1[1480]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2959]),.i2(intermediate_reg_0[2958]),.o(intermediate_reg_1[1479])); 
fsm fsm_inst_1_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2957]),.i2(intermediate_reg_0[2956]),.o(intermediate_reg_1[1478])); 
fsm fsm_inst_1_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2955]),.i2(intermediate_reg_0[2954]),.o(intermediate_reg_1[1477])); 
fsm fsm_inst_1_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2953]),.i2(intermediate_reg_0[2952]),.o(intermediate_reg_1[1476])); 
fsm fsm_inst_1_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2951]),.i2(intermediate_reg_0[2950]),.o(intermediate_reg_1[1475])); 
mux_module mux_module_inst_1_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2949]),.i2(intermediate_reg_0[2948]),.o(intermediate_reg_1[1474]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2947]),.i2(intermediate_reg_0[2946]),.o(intermediate_reg_1[1473])); 
fsm fsm_inst_1_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2945]),.i2(intermediate_reg_0[2944]),.o(intermediate_reg_1[1472])); 
fsm fsm_inst_1_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2943]),.i2(intermediate_reg_0[2942]),.o(intermediate_reg_1[1471])); 
fsm fsm_inst_1_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2941]),.i2(intermediate_reg_0[2940]),.o(intermediate_reg_1[1470])); 
fsm fsm_inst_1_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2939]),.i2(intermediate_reg_0[2938]),.o(intermediate_reg_1[1469])); 
fsm fsm_inst_1_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2937]),.i2(intermediate_reg_0[2936]),.o(intermediate_reg_1[1468])); 
mux_module mux_module_inst_1_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2935]),.i2(intermediate_reg_0[2934]),.o(intermediate_reg_1[1467]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2933]),.i2(intermediate_reg_0[2932]),.o(intermediate_reg_1[1466])); 
fsm fsm_inst_1_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2931]),.i2(intermediate_reg_0[2930]),.o(intermediate_reg_1[1465])); 
mux_module mux_module_inst_1_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2929]),.i2(intermediate_reg_0[2928]),.o(intermediate_reg_1[1464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2927]),.i2(intermediate_reg_0[2926]),.o(intermediate_reg_1[1463]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2925]),.i2(intermediate_reg_0[2924]),.o(intermediate_reg_1[1462])); 
fsm fsm_inst_1_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2923]),.i2(intermediate_reg_0[2922]),.o(intermediate_reg_1[1461])); 
fsm fsm_inst_1_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2921]),.i2(intermediate_reg_0[2920]),.o(intermediate_reg_1[1460])); 
mux_module mux_module_inst_1_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2919]),.i2(intermediate_reg_0[2918]),.o(intermediate_reg_1[1459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2917]),.i2(intermediate_reg_0[2916]),.o(intermediate_reg_1[1458]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2915]),.i2(intermediate_reg_0[2914]),.o(intermediate_reg_1[1457]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2913]),.i2(intermediate_reg_0[2912]),.o(intermediate_reg_1[1456])); 
mux_module mux_module_inst_1_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2911]),.i2(intermediate_reg_0[2910]),.o(intermediate_reg_1[1455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2909]),.i2(intermediate_reg_0[2908]),.o(intermediate_reg_1[1454]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2907]),.i2(intermediate_reg_0[2906]),.o(intermediate_reg_1[1453])); 
mux_module mux_module_inst_1_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2905]),.i2(intermediate_reg_0[2904]),.o(intermediate_reg_1[1452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2903]),.i2(intermediate_reg_0[2902]),.o(intermediate_reg_1[1451]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2901]),.i2(intermediate_reg_0[2900]),.o(intermediate_reg_1[1450])); 
mux_module mux_module_inst_1_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2899]),.i2(intermediate_reg_0[2898]),.o(intermediate_reg_1[1449]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2897]),.i2(intermediate_reg_0[2896]),.o(intermediate_reg_1[1448]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2895]),.i2(intermediate_reg_0[2894]),.o(intermediate_reg_1[1447]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2893]),.i2(intermediate_reg_0[2892]),.o(intermediate_reg_1[1446]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2891]),.i2(intermediate_reg_0[2890]),.o(intermediate_reg_1[1445])); 
mux_module mux_module_inst_1_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2889]),.i2(intermediate_reg_0[2888]),.o(intermediate_reg_1[1444]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2887]),.i2(intermediate_reg_0[2886]),.o(intermediate_reg_1[1443])); 
mux_module mux_module_inst_1_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2885]),.i2(intermediate_reg_0[2884]),.o(intermediate_reg_1[1442]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2883]),.i2(intermediate_reg_0[2882]),.o(intermediate_reg_1[1441]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2881]),.i2(intermediate_reg_0[2880]),.o(intermediate_reg_1[1440])); 
mux_module mux_module_inst_1_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2879]),.i2(intermediate_reg_0[2878]),.o(intermediate_reg_1[1439]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2877]),.i2(intermediate_reg_0[2876]),.o(intermediate_reg_1[1438])); 
mux_module mux_module_inst_1_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2875]),.i2(intermediate_reg_0[2874]),.o(intermediate_reg_1[1437]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2873]),.i2(intermediate_reg_0[2872]),.o(intermediate_reg_1[1436]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2871]),.i2(intermediate_reg_0[2870]),.o(intermediate_reg_1[1435])); 
fsm fsm_inst_1_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2869]),.i2(intermediate_reg_0[2868]),.o(intermediate_reg_1[1434])); 
mux_module mux_module_inst_1_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2867]),.i2(intermediate_reg_0[2866]),.o(intermediate_reg_1[1433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2865]),.i2(intermediate_reg_0[2864]),.o(intermediate_reg_1[1432]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2863]),.i2(intermediate_reg_0[2862]),.o(intermediate_reg_1[1431])); 
fsm fsm_inst_1_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2861]),.i2(intermediate_reg_0[2860]),.o(intermediate_reg_1[1430])); 
fsm fsm_inst_1_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2859]),.i2(intermediate_reg_0[2858]),.o(intermediate_reg_1[1429])); 
fsm fsm_inst_1_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2857]),.i2(intermediate_reg_0[2856]),.o(intermediate_reg_1[1428])); 
mux_module mux_module_inst_1_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2855]),.i2(intermediate_reg_0[2854]),.o(intermediate_reg_1[1427]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2853]),.i2(intermediate_reg_0[2852]),.o(intermediate_reg_1[1426])); 
fsm fsm_inst_1_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2851]),.i2(intermediate_reg_0[2850]),.o(intermediate_reg_1[1425])); 
mux_module mux_module_inst_1_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2849]),.i2(intermediate_reg_0[2848]),.o(intermediate_reg_1[1424]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2847]),.i2(intermediate_reg_0[2846]),.o(intermediate_reg_1[1423])); 
fsm fsm_inst_1_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2845]),.i2(intermediate_reg_0[2844]),.o(intermediate_reg_1[1422])); 
mux_module mux_module_inst_1_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2843]),.i2(intermediate_reg_0[2842]),.o(intermediate_reg_1[1421]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2841]),.i2(intermediate_reg_0[2840]),.o(intermediate_reg_1[1420])); 
fsm fsm_inst_1_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2839]),.i2(intermediate_reg_0[2838]),.o(intermediate_reg_1[1419])); 
mux_module mux_module_inst_1_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2837]),.i2(intermediate_reg_0[2836]),.o(intermediate_reg_1[1418]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2835]),.i2(intermediate_reg_0[2834]),.o(intermediate_reg_1[1417]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2833]),.i2(intermediate_reg_0[2832]),.o(intermediate_reg_1[1416])); 
fsm fsm_inst_1_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2831]),.i2(intermediate_reg_0[2830]),.o(intermediate_reg_1[1415])); 
mux_module mux_module_inst_1_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2829]),.i2(intermediate_reg_0[2828]),.o(intermediate_reg_1[1414]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2827]),.i2(intermediate_reg_0[2826]),.o(intermediate_reg_1[1413]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2825]),.i2(intermediate_reg_0[2824]),.o(intermediate_reg_1[1412])); 
fsm fsm_inst_1_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2823]),.i2(intermediate_reg_0[2822]),.o(intermediate_reg_1[1411])); 
mux_module mux_module_inst_1_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2821]),.i2(intermediate_reg_0[2820]),.o(intermediate_reg_1[1410]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2819]),.i2(intermediate_reg_0[2818]),.o(intermediate_reg_1[1409]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2817]),.i2(intermediate_reg_0[2816]),.o(intermediate_reg_1[1408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2815]),.i2(intermediate_reg_0[2814]),.o(intermediate_reg_1[1407]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2813]),.i2(intermediate_reg_0[2812]),.o(intermediate_reg_1[1406]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2811]),.i2(intermediate_reg_0[2810]),.o(intermediate_reg_1[1405])); 
mux_module mux_module_inst_1_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2809]),.i2(intermediate_reg_0[2808]),.o(intermediate_reg_1[1404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2807]),.i2(intermediate_reg_0[2806]),.o(intermediate_reg_1[1403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2805]),.i2(intermediate_reg_0[2804]),.o(intermediate_reg_1[1402]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2803]),.i2(intermediate_reg_0[2802]),.o(intermediate_reg_1[1401])); 
fsm fsm_inst_1_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2801]),.i2(intermediate_reg_0[2800]),.o(intermediate_reg_1[1400])); 
mux_module mux_module_inst_1_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2799]),.i2(intermediate_reg_0[2798]),.o(intermediate_reg_1[1399]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2797]),.i2(intermediate_reg_0[2796]),.o(intermediate_reg_1[1398])); 
fsm fsm_inst_1_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2795]),.i2(intermediate_reg_0[2794]),.o(intermediate_reg_1[1397])); 
fsm fsm_inst_1_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2793]),.i2(intermediate_reg_0[2792]),.o(intermediate_reg_1[1396])); 
mux_module mux_module_inst_1_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2791]),.i2(intermediate_reg_0[2790]),.o(intermediate_reg_1[1395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2789]),.i2(intermediate_reg_0[2788]),.o(intermediate_reg_1[1394]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2787]),.i2(intermediate_reg_0[2786]),.o(intermediate_reg_1[1393])); 
fsm fsm_inst_1_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2785]),.i2(intermediate_reg_0[2784]),.o(intermediate_reg_1[1392])); 
fsm fsm_inst_1_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2783]),.i2(intermediate_reg_0[2782]),.o(intermediate_reg_1[1391])); 
mux_module mux_module_inst_1_1649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2781]),.i2(intermediate_reg_0[2780]),.o(intermediate_reg_1[1390]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2779]),.i2(intermediate_reg_0[2778]),.o(intermediate_reg_1[1389]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2777]),.i2(intermediate_reg_0[2776]),.o(intermediate_reg_1[1388]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2775]),.i2(intermediate_reg_0[2774]),.o(intermediate_reg_1[1387]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2773]),.i2(intermediate_reg_0[2772]),.o(intermediate_reg_1[1386])); 
fsm fsm_inst_1_1654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2771]),.i2(intermediate_reg_0[2770]),.o(intermediate_reg_1[1385])); 
mux_module mux_module_inst_1_1655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2769]),.i2(intermediate_reg_0[2768]),.o(intermediate_reg_1[1384]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2767]),.i2(intermediate_reg_0[2766]),.o(intermediate_reg_1[1383]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2765]),.i2(intermediate_reg_0[2764]),.o(intermediate_reg_1[1382])); 
fsm fsm_inst_1_1658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2763]),.i2(intermediate_reg_0[2762]),.o(intermediate_reg_1[1381])); 
mux_module mux_module_inst_1_1659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2761]),.i2(intermediate_reg_0[2760]),.o(intermediate_reg_1[1380]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2759]),.i2(intermediate_reg_0[2758]),.o(intermediate_reg_1[1379])); 
mux_module mux_module_inst_1_1661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2757]),.i2(intermediate_reg_0[2756]),.o(intermediate_reg_1[1378]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2755]),.i2(intermediate_reg_0[2754]),.o(intermediate_reg_1[1377]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2753]),.i2(intermediate_reg_0[2752]),.o(intermediate_reg_1[1376])); 
mux_module mux_module_inst_1_1664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2751]),.i2(intermediate_reg_0[2750]),.o(intermediate_reg_1[1375]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2749]),.i2(intermediate_reg_0[2748]),.o(intermediate_reg_1[1374])); 
mux_module mux_module_inst_1_1666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2747]),.i2(intermediate_reg_0[2746]),.o(intermediate_reg_1[1373]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2745]),.i2(intermediate_reg_0[2744]),.o(intermediate_reg_1[1372])); 
mux_module mux_module_inst_1_1668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2743]),.i2(intermediate_reg_0[2742]),.o(intermediate_reg_1[1371]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2741]),.i2(intermediate_reg_0[2740]),.o(intermediate_reg_1[1370])); 
fsm fsm_inst_1_1670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2739]),.i2(intermediate_reg_0[2738]),.o(intermediate_reg_1[1369])); 
mux_module mux_module_inst_1_1671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2737]),.i2(intermediate_reg_0[2736]),.o(intermediate_reg_1[1368]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2735]),.i2(intermediate_reg_0[2734]),.o(intermediate_reg_1[1367]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2733]),.i2(intermediate_reg_0[2732]),.o(intermediate_reg_1[1366]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2731]),.i2(intermediate_reg_0[2730]),.o(intermediate_reg_1[1365])); 
fsm fsm_inst_1_1675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2729]),.i2(intermediate_reg_0[2728]),.o(intermediate_reg_1[1364])); 
mux_module mux_module_inst_1_1676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2727]),.i2(intermediate_reg_0[2726]),.o(intermediate_reg_1[1363]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2725]),.i2(intermediate_reg_0[2724]),.o(intermediate_reg_1[1362]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2723]),.i2(intermediate_reg_0[2722]),.o(intermediate_reg_1[1361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2721]),.i2(intermediate_reg_0[2720]),.o(intermediate_reg_1[1360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2719]),.i2(intermediate_reg_0[2718]),.o(intermediate_reg_1[1359]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2717]),.i2(intermediate_reg_0[2716]),.o(intermediate_reg_1[1358])); 
mux_module mux_module_inst_1_1682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2715]),.i2(intermediate_reg_0[2714]),.o(intermediate_reg_1[1357]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2713]),.i2(intermediate_reg_0[2712]),.o(intermediate_reg_1[1356])); 
mux_module mux_module_inst_1_1684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2711]),.i2(intermediate_reg_0[2710]),.o(intermediate_reg_1[1355]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2709]),.i2(intermediate_reg_0[2708]),.o(intermediate_reg_1[1354])); 
fsm fsm_inst_1_1686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2707]),.i2(intermediate_reg_0[2706]),.o(intermediate_reg_1[1353])); 
fsm fsm_inst_1_1687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2705]),.i2(intermediate_reg_0[2704]),.o(intermediate_reg_1[1352])); 
fsm fsm_inst_1_1688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2703]),.i2(intermediate_reg_0[2702]),.o(intermediate_reg_1[1351])); 
fsm fsm_inst_1_1689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2701]),.i2(intermediate_reg_0[2700]),.o(intermediate_reg_1[1350])); 
fsm fsm_inst_1_1690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2699]),.i2(intermediate_reg_0[2698]),.o(intermediate_reg_1[1349])); 
fsm fsm_inst_1_1691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2697]),.i2(intermediate_reg_0[2696]),.o(intermediate_reg_1[1348])); 
fsm fsm_inst_1_1692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2695]),.i2(intermediate_reg_0[2694]),.o(intermediate_reg_1[1347])); 
mux_module mux_module_inst_1_1693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2693]),.i2(intermediate_reg_0[2692]),.o(intermediate_reg_1[1346]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2691]),.i2(intermediate_reg_0[2690]),.o(intermediate_reg_1[1345])); 
fsm fsm_inst_1_1695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2689]),.i2(intermediate_reg_0[2688]),.o(intermediate_reg_1[1344])); 
mux_module mux_module_inst_1_1696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339])); 
fsm fsm_inst_1_1701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338])); 
mux_module mux_module_inst_1_1702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335])); 
mux_module mux_module_inst_1_1705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330])); 
mux_module mux_module_inst_1_1710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328])); 
mux_module mux_module_inst_1_1712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326])); 
mux_module mux_module_inst_1_1714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324])); 
mux_module mux_module_inst_1_1716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322])); 
mux_module mux_module_inst_1_1718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320])); 
mux_module mux_module_inst_1_1720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317])); 
mux_module mux_module_inst_1_1723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315])); 
mux_module mux_module_inst_1_1725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313])); 
mux_module mux_module_inst_1_1727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309])); 
fsm fsm_inst_1_1731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308])); 
fsm fsm_inst_1_1732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307])); 
mux_module mux_module_inst_1_1733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305])); 
fsm fsm_inst_1_1735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304])); 
fsm fsm_inst_1_1736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303])); 
mux_module mux_module_inst_1_1737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298])); 
fsm fsm_inst_1_1742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297])); 
fsm fsm_inst_1_1743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296])); 
fsm fsm_inst_1_1744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295])); 
fsm fsm_inst_1_1745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294])); 
mux_module mux_module_inst_1_1746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291])); 
fsm fsm_inst_1_1749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290])); 
mux_module mux_module_inst_1_1750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286])); 
mux_module mux_module_inst_1_1754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284])); 
mux_module mux_module_inst_1_1756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282])); 
mux_module mux_module_inst_1_1758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280])); 
mux_module mux_module_inst_1_1760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277])); 
mux_module mux_module_inst_1_1763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275])); 
mux_module mux_module_inst_1_1765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273])); 
fsm fsm_inst_1_1767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272])); 
fsm fsm_inst_1_1768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271])); 
fsm fsm_inst_1_1769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270])); 
fsm fsm_inst_1_1770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269])); 
fsm fsm_inst_1_1771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268])); 
mux_module mux_module_inst_1_1772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266])); 
mux_module mux_module_inst_1_1774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258])); 
fsm fsm_inst_1_1782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257])); 
mux_module mux_module_inst_1_1783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254])); 
fsm fsm_inst_1_1786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253])); 
fsm fsm_inst_1_1787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252])); 
mux_module mux_module_inst_1_1788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250])); 
mux_module mux_module_inst_1_1790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248])); 
mux_module mux_module_inst_1_1792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246])); 
fsm fsm_inst_1_1794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245])); 
fsm fsm_inst_1_1795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244])); 
fsm fsm_inst_1_1796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243])); 
mux_module mux_module_inst_1_1797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
fsm fsm_inst_1_1800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239])); 
fsm fsm_inst_1_1801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238])); 
mux_module mux_module_inst_1_1802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234])); 
mux_module mux_module_inst_1_1806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230])); 
fsm fsm_inst_1_1810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229])); 
fsm fsm_inst_1_1811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228])); 
mux_module mux_module_inst_1_1812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
fsm fsm_inst_1_1814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225])); 
mux_module mux_module_inst_1_1815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223])); 
fsm fsm_inst_1_1817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222])); 
fsm fsm_inst_1_1818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
mux_module mux_module_inst_1_1819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219])); 
mux_module mux_module_inst_1_1821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216])); 
fsm fsm_inst_1_1824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215])); 
mux_module mux_module_inst_1_1825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213])); 
mux_module mux_module_inst_1_1827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211])); 
fsm fsm_inst_1_1829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210])); 
fsm fsm_inst_1_1830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209])); 
fsm fsm_inst_1_1831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208])); 
fsm fsm_inst_1_1832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207])); 
fsm fsm_inst_1_1833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206])); 
fsm fsm_inst_1_1834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205])); 
fsm fsm_inst_1_1835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204])); 
mux_module mux_module_inst_1_1836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201])); 
fsm fsm_inst_1_1839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200])); 
mux_module mux_module_inst_1_1840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197])); 
mux_module mux_module_inst_1_1843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188])); 
mux_module mux_module_inst_1_1852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185])); 
fsm fsm_inst_1_1855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184])); 
mux_module mux_module_inst_1_1856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181])); 
mux_module mux_module_inst_1_1859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179])); 
mux_module mux_module_inst_1_1861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176])); 
fsm fsm_inst_1_1864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175])); 
fsm fsm_inst_1_1865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174])); 
mux_module mux_module_inst_1_1866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172])); 
fsm fsm_inst_1_1868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171])); 
fsm fsm_inst_1_1869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170])); 
mux_module mux_module_inst_1_1870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167])); 
fsm fsm_inst_1_1873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166])); 
mux_module mux_module_inst_1_1874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164])); 
mux_module mux_module_inst_1_1876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
fsm fsm_inst_1_1883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156])); 
fsm fsm_inst_1_1884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155])); 
fsm fsm_inst_1_1885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154])); 
fsm fsm_inst_1_1886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153])); 
mux_module mux_module_inst_1_1887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151])); 
fsm fsm_inst_1_1889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150])); 
fsm fsm_inst_1_1890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149])); 
fsm fsm_inst_1_1891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
fsm fsm_inst_1_1892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147])); 
mux_module mux_module_inst_1_1893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143])); 
mux_module mux_module_inst_1_1897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141])); 
mux_module mux_module_inst_1_1899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138])); 
mux_module mux_module_inst_1_1902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136])); 
mux_module mux_module_inst_1_1904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
fsm fsm_inst_1_1910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129])); 
fsm fsm_inst_1_1911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128])); 
mux_module mux_module_inst_1_1912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126])); 
mux_module mux_module_inst_1_1914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121])); 
fsm fsm_inst_1_1919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120])); 
fsm fsm_inst_1_1920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
mux_module mux_module_inst_1_1921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116])); 
mux_module mux_module_inst_1_1924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114])); 
fsm fsm_inst_1_1926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113])); 
mux_module mux_module_inst_1_1927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110])); 
mux_module mux_module_inst_1_1930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107])); 
fsm fsm_inst_1_1933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106])); 
fsm fsm_inst_1_1934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
mux_module mux_module_inst_1_1935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
mux_module mux_module_inst_1_1937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
mux_module mux_module_inst_1_1939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
fsm fsm_inst_1_1947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
fsm fsm_inst_1_1948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
mux_module mux_module_inst_1_1949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
mux_module mux_module_inst_1_1951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
fsm fsm_inst_1_1953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086])); 
fsm fsm_inst_1_1954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085])); 
fsm fsm_inst_1_1955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084])); 
fsm fsm_inst_1_1956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
mux_module mux_module_inst_1_1957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081])); 
mux_module mux_module_inst_1_1959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079])); 
mux_module mux_module_inst_1_1961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077])); 
mux_module mux_module_inst_1_1963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075])); 
fsm fsm_inst_1_1965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074])); 
fsm fsm_inst_1_1966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
mux_module mux_module_inst_1_1967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071])); 
fsm fsm_inst_1_1969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070])); 
fsm fsm_inst_1_1970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069])); 
mux_module mux_module_inst_1_1971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066])); 
mux_module mux_module_inst_1_1974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064])); 
fsm fsm_inst_1_1976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063])); 
fsm fsm_inst_1_1977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062])); 
fsm fsm_inst_1_1978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061])); 
mux_module mux_module_inst_1_1979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059])); 
mux_module mux_module_inst_1_1981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055])); 
fsm fsm_inst_1_1985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054])); 
fsm fsm_inst_1_1986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053])); 
mux_module mux_module_inst_1_1987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051])); 
mux_module mux_module_inst_1_1989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049])); 
mux_module mux_module_inst_1_1991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
mux_module mux_module_inst_1_1993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
mux_module mux_module_inst_1_1998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040])); 
fsm fsm_inst_1_2000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039])); 
mux_module mux_module_inst_1_2001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036])); 
mux_module mux_module_inst_1_2004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
mux_module mux_module_inst_1_2009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029])); 
fsm fsm_inst_1_2011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
mux_module mux_module_inst_1_2012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
mux_module mux_module_inst_1_2015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
fsm fsm_inst_1_2017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022])); 
mux_module mux_module_inst_1_2018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
fsm fsm_inst_1_2021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018])); 
fsm fsm_inst_1_2022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017])); 
fsm fsm_inst_1_2023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016])); 
mux_module mux_module_inst_1_2024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
fsm fsm_inst_1_2026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013])); 
fsm fsm_inst_1_2027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012])); 
fsm fsm_inst_1_2028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011])); 
mux_module mux_module_inst_1_2029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009])); 
fsm fsm_inst_1_2031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
fsm fsm_inst_1_2032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
fsm fsm_inst_1_2033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006])); 
fsm fsm_inst_1_2034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
mux_module mux_module_inst_1_2035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001])); 
fsm fsm_inst_1_2039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
mux_module mux_module_inst_1_2040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
mux_module mux_module_inst_1_2042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
fsm fsm_inst_1_2045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
fsm fsm_inst_1_2046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
fsm fsm_inst_1_2047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
mux_module mux_module_inst_1_2048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
fsm fsm_inst_1_2050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
mux_module mux_module_inst_1_2051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
mux_module mux_module_inst_1_2053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
mux_module mux_module_inst_1_2058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
mux_module mux_module_inst_1_2064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973])); 
fsm fsm_inst_1_2067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
fsm fsm_inst_1_2068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971])); 
mux_module mux_module_inst_1_2069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
fsm fsm_inst_1_2071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
fsm fsm_inst_1_2072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
mux_module mux_module_inst_1_2073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
mux_module mux_module_inst_1_2076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
fsm fsm_inst_1_2079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
mux_module mux_module_inst_1_2080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
mux_module mux_module_inst_1_2082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
fsm fsm_inst_1_2084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
mux_module mux_module_inst_1_2085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
mux_module mux_module_inst_1_2087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950])); 
fsm fsm_inst_1_2090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
mux_module mux_module_inst_1_2091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
mux_module mux_module_inst_1_2093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
fsm fsm_inst_1_2098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
mux_module mux_module_inst_1_2099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
fsm fsm_inst_1_2101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
mux_module mux_module_inst_1_2102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
mux_module mux_module_inst_1_2104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
fsm fsm_inst_1_2106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
mux_module mux_module_inst_1_2107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
fsm fsm_inst_1_2111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
mux_module mux_module_inst_1_2112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
fsm fsm_inst_1_2114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
mux_module mux_module_inst_1_2115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
fsm fsm_inst_1_2117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
fsm fsm_inst_1_2118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
fsm fsm_inst_1_2119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
fsm fsm_inst_1_2120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
fsm fsm_inst_1_2121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
mux_module mux_module_inst_1_2122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
mux_module mux_module_inst_1_2124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
fsm fsm_inst_1_2127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
mux_module mux_module_inst_1_2128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
fsm fsm_inst_1_2130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
fsm fsm_inst_1_2131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
mux_module mux_module_inst_1_2132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906])); 
mux_module mux_module_inst_1_2134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
mux_module mux_module_inst_1_2136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
fsm fsm_inst_1_2138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
fsm fsm_inst_1_2139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
fsm fsm_inst_1_2140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
fsm fsm_inst_1_2141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
mux_module mux_module_inst_1_2142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
mux_module mux_module_inst_1_2144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
mux_module mux_module_inst_1_2146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
fsm fsm_inst_1_2148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
mux_module mux_module_inst_1_2149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
fsm fsm_inst_1_2151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
fsm fsm_inst_1_2152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
mux_module mux_module_inst_1_2153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
fsm fsm_inst_1_2157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
fsm fsm_inst_1_2158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
fsm fsm_inst_1_2159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
mux_module mux_module_inst_1_2160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
fsm fsm_inst_1_2163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
mux_module mux_module_inst_1_2164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
fsm fsm_inst_1_2167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
fsm fsm_inst_1_2168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
fsm fsm_inst_1_2169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
mux_module mux_module_inst_1_2170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
fsm fsm_inst_1_2172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
mux_module mux_module_inst_1_2173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
fsm fsm_inst_1_2177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862])); 
mux_module mux_module_inst_1_2178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
fsm fsm_inst_1_2180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859])); 
fsm fsm_inst_1_2181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
mux_module mux_module_inst_1_2182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
mux_module mux_module_inst_1_2187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
fsm fsm_inst_1_2189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
mux_module mux_module_inst_1_2190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
mux_module mux_module_inst_1_2195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
mux_module mux_module_inst_1_2197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
fsm fsm_inst_1_2200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
mux_module mux_module_inst_1_2201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
fsm fsm_inst_1_2204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
mux_module mux_module_inst_1_2205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832])); 
mux_module mux_module_inst_1_2208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
mux_module mux_module_inst_1_2212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
fsm fsm_inst_1_2218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
mux_module mux_module_inst_1_2219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
fsm fsm_inst_1_2225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
fsm fsm_inst_1_2226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
fsm fsm_inst_1_2227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
fsm fsm_inst_1_2228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
mux_module mux_module_inst_1_2229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
mux_module mux_module_inst_1_2232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
mux_module mux_module_inst_1_2235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803])); 
mux_module mux_module_inst_1_2237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
mux_module mux_module_inst_1_2239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
fsm fsm_inst_1_2241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
fsm fsm_inst_1_2242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
fsm fsm_inst_1_2243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
mux_module mux_module_inst_1_2244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
fsm fsm_inst_1_2247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
fsm fsm_inst_1_2248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
mux_module mux_module_inst_1_2249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
mux_module mux_module_inst_1_2251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
fsm fsm_inst_1_2254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
fsm fsm_inst_1_2255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784])); 
mux_module mux_module_inst_1_2256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
fsm fsm_inst_1_2258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
mux_module mux_module_inst_1_2259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
fsm fsm_inst_1_2262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
fsm fsm_inst_1_2263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
mux_module mux_module_inst_1_2264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
mux_module mux_module_inst_1_2266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
mux_module mux_module_inst_1_2268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
mux_module mux_module_inst_1_2273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
mux_module mux_module_inst_1_2278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
fsm fsm_inst_1_2283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
mux_module mux_module_inst_1_2284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
mux_module mux_module_inst_1_2286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
mux_module mux_module_inst_1_2289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
mux_module mux_module_inst_1_2292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
mux_module mux_module_inst_1_2294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
mux_module mux_module_inst_1_2296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
fsm fsm_inst_1_2299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
fsm fsm_inst_1_2300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
mux_module mux_module_inst_1_2301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
fsm fsm_inst_1_2303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
mux_module mux_module_inst_1_2304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
fsm fsm_inst_1_2306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
fsm fsm_inst_1_2307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
mux_module mux_module_inst_1_2308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
mux_module mux_module_inst_1_2311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
mux_module mux_module_inst_1_2316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
fsm fsm_inst_1_2319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
mux_module mux_module_inst_1_2320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
fsm fsm_inst_1_2323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
mux_module mux_module_inst_1_2324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
mux_module mux_module_inst_1_2326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
fsm fsm_inst_1_2329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
fsm fsm_inst_1_2330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
fsm fsm_inst_1_2331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
mux_module mux_module_inst_1_2332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
fsm fsm_inst_1_2335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
mux_module mux_module_inst_1_2336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
mux_module mux_module_inst_1_2340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
fsm fsm_inst_1_2346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
mux_module mux_module_inst_1_2347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
mux_module mux_module_inst_1_2352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
fsm fsm_inst_1_2355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
mux_module mux_module_inst_1_2356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
fsm fsm_inst_1_2358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
fsm fsm_inst_1_2359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
fsm fsm_inst_1_2360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
mux_module mux_module_inst_1_2361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
mux_module mux_module_inst_1_2364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
fsm fsm_inst_1_2368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
fsm fsm_inst_1_2369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
mux_module mux_module_inst_1_2370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
fsm fsm_inst_1_2375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
mux_module mux_module_inst_1_2376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
mux_module mux_module_inst_1_2378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
fsm fsm_inst_1_2380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_2381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
fsm fsm_inst_1_2382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
mux_module mux_module_inst_1_2383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
fsm fsm_inst_1_2386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
mux_module mux_module_inst_1_2387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
fsm fsm_inst_1_2391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
mux_module mux_module_inst_1_2392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
fsm fsm_inst_1_2395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
fsm fsm_inst_1_2396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
mux_module mux_module_inst_1_2397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640])); 
mux_module mux_module_inst_1_2400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
mux_module mux_module_inst_1_2402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
fsm fsm_inst_1_2406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
mux_module mux_module_inst_1_2407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
mux_module mux_module_inst_1_2409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
fsm fsm_inst_1_2411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
mux_module mux_module_inst_1_2412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626])); 
fsm fsm_inst_1_2414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
fsm fsm_inst_1_2415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
fsm fsm_inst_1_2416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
fsm fsm_inst_1_2417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
mux_module mux_module_inst_1_2418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
fsm fsm_inst_1_2424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
fsm fsm_inst_1_2425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
mux_module mux_module_inst_1_2426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
fsm fsm_inst_1_2428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
mux_module mux_module_inst_1_2429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
fsm fsm_inst_1_2432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
fsm fsm_inst_1_2433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
mux_module mux_module_inst_1_2434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
fsm fsm_inst_1_2436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
mux_module mux_module_inst_1_2437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
fsm fsm_inst_1_2439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
mux_module mux_module_inst_1_2440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
fsm fsm_inst_1_2443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
mux_module mux_module_inst_1_2444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_2446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
fsm fsm_inst_1_2447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
mux_module mux_module_inst_1_2448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
mux_module mux_module_inst_1_2450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
mux_module mux_module_inst_1_2452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
mux_module mux_module_inst_1_2454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
mux_module mux_module_inst_1_2456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
mux_module mux_module_inst_1_2458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
mux_module mux_module_inst_1_2460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
fsm fsm_inst_1_2462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
fsm fsm_inst_1_2463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
fsm fsm_inst_1_2464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
fsm fsm_inst_1_2465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
mux_module mux_module_inst_1_2466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
fsm fsm_inst_1_2469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
fsm fsm_inst_1_2470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
fsm fsm_inst_1_2471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
mux_module mux_module_inst_1_2472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565])); 
fsm fsm_inst_1_2475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
fsm fsm_inst_1_2476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
mux_module mux_module_inst_1_2477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
fsm fsm_inst_1_2480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
mux_module mux_module_inst_1_2481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
fsm fsm_inst_1_2485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
fsm fsm_inst_1_2486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_2487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
mux_module mux_module_inst_1_2488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
mux_module mux_module_inst_1_2490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
fsm fsm_inst_1_2493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
mux_module mux_module_inst_1_2494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
fsm fsm_inst_1_2496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
fsm fsm_inst_1_2497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
fsm fsm_inst_1_2498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
mux_module mux_module_inst_1_2499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
mux_module mux_module_inst_1_2503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_2505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
mux_module mux_module_inst_1_2506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
fsm fsm_inst_1_2509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
mux_module mux_module_inst_1_2510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
mux_module mux_module_inst_1_2513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
fsm fsm_inst_1_2515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
mux_module mux_module_inst_1_2516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
fsm fsm_inst_1_2519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
fsm fsm_inst_1_2520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
mux_module mux_module_inst_1_2521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
mux_module mux_module_inst_1_2523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
fsm fsm_inst_1_2525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
fsm fsm_inst_1_2526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
fsm fsm_inst_1_2527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
fsm fsm_inst_1_2528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
mux_module mux_module_inst_1_2529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508])); 
fsm fsm_inst_1_2532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
mux_module mux_module_inst_1_2533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
mux_module mux_module_inst_1_2535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
mux_module mux_module_inst_1_2537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
mux_module mux_module_inst_1_2539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
mux_module mux_module_inst_1_2541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
mux_module mux_module_inst_1_2543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
fsm fsm_inst_1_2546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
mux_module mux_module_inst_1_2547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
mux_module mux_module_inst_1_2549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
fsm fsm_inst_1_2552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
fsm fsm_inst_1_2553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
mux_module mux_module_inst_1_2554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
fsm fsm_inst_1_2557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_2558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
mux_module mux_module_inst_1_2561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_2563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
mux_module mux_module_inst_1_2564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
fsm fsm_inst_1_2566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
fsm fsm_inst_1_2567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
mux_module mux_module_inst_1_2568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
fsm fsm_inst_1_2570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
fsm fsm_inst_1_2571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
mux_module mux_module_inst_1_2572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
mux_module mux_module_inst_1_2574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
fsm fsm_inst_1_2581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
mux_module mux_module_inst_1_2582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
mux_module mux_module_inst_1_2584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
fsm fsm_inst_1_2586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
fsm fsm_inst_1_2587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
fsm fsm_inst_1_2588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
fsm fsm_inst_1_2589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
mux_module mux_module_inst_1_2590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
fsm fsm_inst_1_2592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
fsm fsm_inst_1_2593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
mux_module mux_module_inst_1_2594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
mux_module mux_module_inst_1_2596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
mux_module mux_module_inst_1_2598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
fsm fsm_inst_1_2600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
fsm fsm_inst_1_2601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
fsm fsm_inst_1_2602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
mux_module mux_module_inst_1_2603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
mux_module mux_module_inst_1_2607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
fsm fsm_inst_1_2609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
mux_module mux_module_inst_1_2610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
mux_module mux_module_inst_1_2620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
fsm fsm_inst_1_2625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
fsm fsm_inst_1_2626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
fsm fsm_inst_1_2627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
fsm fsm_inst_1_2628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
mux_module mux_module_inst_1_2629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
fsm fsm_inst_1_2631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
mux_module mux_module_inst_1_2632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
fsm fsm_inst_1_2634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405])); 
mux_module mux_module_inst_1_2635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
mux_module mux_module_inst_1_2637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
mux_module mux_module_inst_1_2639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
fsm fsm_inst_1_2643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
fsm fsm_inst_1_2644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
fsm fsm_inst_1_2645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_2646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_2647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
fsm fsm_inst_1_2649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
fsm fsm_inst_1_2650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
mux_module mux_module_inst_1_2651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
fsm fsm_inst_1_2654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_2655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
mux_module mux_module_inst_1_2658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
fsm fsm_inst_1_2660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
fsm fsm_inst_1_2661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
fsm fsm_inst_1_2662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_2663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
fsm fsm_inst_1_2664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
fsm fsm_inst_1_2665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
fsm fsm_inst_1_2666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
fsm fsm_inst_1_2667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
fsm fsm_inst_1_2668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
mux_module mux_module_inst_1_2669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
mux_module mux_module_inst_1_2672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
mux_module mux_module_inst_1_2674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
mux_module mux_module_inst_1_2676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
mux_module mux_module_inst_1_2678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
fsm fsm_inst_1_2682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
fsm fsm_inst_1_2683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
mux_module mux_module_inst_1_2684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
fsm fsm_inst_1_2686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
mux_module mux_module_inst_1_2687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
fsm fsm_inst_1_2691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
mux_module mux_module_inst_1_2692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
fsm fsm_inst_1_2694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
fsm fsm_inst_1_2695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
fsm fsm_inst_1_2696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
fsm fsm_inst_1_2697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
fsm fsm_inst_1_2698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
mux_module mux_module_inst_1_2699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
fsm fsm_inst_1_2701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
mux_module mux_module_inst_1_2702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
mux_module mux_module_inst_1_2705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
fsm fsm_inst_1_2709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330])); 
mux_module mux_module_inst_1_2710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
fsm fsm_inst_1_2713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
fsm fsm_inst_1_2714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
mux_module mux_module_inst_1_2715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
fsm fsm_inst_1_2720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
mux_module mux_module_inst_1_2721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
mux_module mux_module_inst_1_2731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
mux_module mux_module_inst_1_2735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
mux_module mux_module_inst_1_2740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
mux_module mux_module_inst_1_2744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
mux_module mux_module_inst_1_2746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
fsm fsm_inst_1_2749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
fsm fsm_inst_1_2750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
mux_module mux_module_inst_1_2751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284])); 
mux_module mux_module_inst_1_2756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
mux_module mux_module_inst_1_2762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
fsm fsm_inst_1_2765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
fsm fsm_inst_1_2766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
mux_module mux_module_inst_1_2767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
mux_module mux_module_inst_1_2772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
fsm fsm_inst_1_2775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
mux_module mux_module_inst_1_2776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_2779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
fsm fsm_inst_1_2780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
fsm fsm_inst_1_2781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
fsm fsm_inst_1_2782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
fsm fsm_inst_1_2783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
fsm fsm_inst_1_2784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
mux_module mux_module_inst_1_2785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
fsm fsm_inst_1_2788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
fsm fsm_inst_1_2789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
mux_module mux_module_inst_1_2790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
mux_module mux_module_inst_1_2792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
mux_module mux_module_inst_1_2794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
fsm fsm_inst_1_2797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
fsm fsm_inst_1_2798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
fsm fsm_inst_1_2799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
fsm fsm_inst_1_2800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239])); 
fsm fsm_inst_1_2801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
mux_module mux_module_inst_1_2802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
mux_module mux_module_inst_1_2804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
mux_module mux_module_inst_1_2807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
fsm fsm_inst_1_2810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
fsm fsm_inst_1_2811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
fsm fsm_inst_1_2812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
mux_module mux_module_inst_1_2813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
mux_module mux_module_inst_1_2816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
fsm fsm_inst_1_2818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
fsm fsm_inst_1_2819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
fsm fsm_inst_1_2820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
fsm fsm_inst_1_2821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
fsm fsm_inst_1_2822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
mux_module mux_module_inst_1_2823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
fsm fsm_inst_1_2825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
fsm fsm_inst_1_2826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
fsm fsm_inst_1_2827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
fsm fsm_inst_1_2828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
fsm fsm_inst_1_2829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
fsm fsm_inst_1_2830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
fsm fsm_inst_1_2831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
mux_module mux_module_inst_1_2832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
fsm fsm_inst_1_2835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
fsm fsm_inst_1_2836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
fsm fsm_inst_1_2837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
mux_module mux_module_inst_1_2838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
fsm fsm_inst_1_2841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
fsm fsm_inst_1_2842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
fsm fsm_inst_1_2843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
fsm fsm_inst_1_2844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
mux_module mux_module_inst_1_2845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
fsm fsm_inst_1_2848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191])); 
fsm fsm_inst_1_2849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
mux_module mux_module_inst_1_2850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
fsm fsm_inst_1_2852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
fsm fsm_inst_1_2853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
fsm fsm_inst_1_2854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
fsm fsm_inst_1_2855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
fsm fsm_inst_1_2856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
fsm fsm_inst_1_2857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
mux_module mux_module_inst_1_2858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
fsm fsm_inst_1_2860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
fsm fsm_inst_1_2861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
fsm fsm_inst_1_2862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
fsm fsm_inst_1_2863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
mux_module mux_module_inst_1_2864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
fsm fsm_inst_1_2867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
mux_module mux_module_inst_1_2868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169])); 
fsm fsm_inst_1_2871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
mux_module mux_module_inst_1_2872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
fsm fsm_inst_1_2874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
mux_module mux_module_inst_1_2875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161])); 
fsm fsm_inst_1_2879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
fsm fsm_inst_1_2880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
mux_module mux_module_inst_1_2881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
fsm fsm_inst_1_2883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
fsm fsm_inst_1_2884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
mux_module mux_module_inst_1_2885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
fsm fsm_inst_1_2888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
mux_module mux_module_inst_1_2889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
fsm fsm_inst_1_2891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
fsm fsm_inst_1_2892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
mux_module mux_module_inst_1_2893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
fsm fsm_inst_1_2895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
mux_module mux_module_inst_1_2896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_2898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
fsm fsm_inst_1_2899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
fsm fsm_inst_1_2900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
fsm fsm_inst_1_2901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
fsm fsm_inst_1_2902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
mux_module mux_module_inst_1_2903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
mux_module mux_module_inst_1_2907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
mux_module mux_module_inst_1_2909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
mux_module mux_module_inst_1_2911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
fsm fsm_inst_1_2913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
fsm fsm_inst_1_2914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
mux_module mux_module_inst_1_2915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
fsm fsm_inst_1_2917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
mux_module mux_module_inst_1_2918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
mux_module mux_module_inst_1_2920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
mux_module mux_module_inst_1_2922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
mux_module mux_module_inst_1_2924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
fsm fsm_inst_1_2927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
mux_module mux_module_inst_1_2928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
mux_module mux_module_inst_1_2930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
fsm fsm_inst_1_2933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
mux_module mux_module_inst_1_2934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
mux_module mux_module_inst_1_2936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
mux_module mux_module_inst_1_2938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
mux_module mux_module_inst_1_2942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
mux_module mux_module_inst_1_2944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
fsm fsm_inst_1_2947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
mux_module mux_module_inst_1_2948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
fsm fsm_inst_1_2950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89])); 
fsm fsm_inst_1_2951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
fsm fsm_inst_1_2952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
fsm fsm_inst_1_2953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
mux_module mux_module_inst_1_2954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
fsm fsm_inst_1_2956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
mux_module mux_module_inst_1_2957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
mux_module mux_module_inst_1_2959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
fsm fsm_inst_1_2962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
mux_module mux_module_inst_1_2963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
fsm fsm_inst_1_2967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
fsm fsm_inst_1_2968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
fsm fsm_inst_1_2969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_2970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
mux_module mux_module_inst_1_2972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_2974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
fsm fsm_inst_1_2977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
mux_module mux_module_inst_1_2978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
mux_module mux_module_inst_1_2980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
fsm fsm_inst_1_2984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
fsm fsm_inst_1_2985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
fsm fsm_inst_1_2986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53])); 
fsm fsm_inst_1_2987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
fsm fsm_inst_1_2988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
fsm fsm_inst_1_2989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_2990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
mux_module mux_module_inst_1_2991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
mux_module mux_module_inst_1_2994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
fsm fsm_inst_1_2998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_2999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
fsm fsm_inst_1_3002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
mux_module mux_module_inst_1_3003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_3005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
mux_module mux_module_inst_1_3006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
mux_module mux_module_inst_1_3009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
fsm fsm_inst_1_3012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
mux_module mux_module_inst_1_3013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
fsm fsm_inst_1_3016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
fsm fsm_inst_1_3017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
fsm fsm_inst_1_3018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
mux_module mux_module_inst_1_3019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
mux_module mux_module_inst_1_3027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
mux_module mux_module_inst_1_3030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
mux_module mux_module_inst_1_3032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_3035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
mux_module mux_module_inst_1_3036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
fsm fsm_inst_1_3038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
mux_module mux_module_inst_1_3039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
always@(posedge clk) begin 
outp [3039:0] <= intermediate_reg_1; 
outp[4991:3040] <= intermediate_reg_1[1951:0] ; 
end 
endmodule 
 

module interface_21(input reg [831:0] inp, output reg [2063:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[831:0] <= inp ; 
outp[1663:832] <= inp ; 
outp[2063:1664] <= inp[399:0] ; 
end 
endmodule 

module interface_22(input reg [2055:0] inp, output reg [311:0] outp, input clk, input reset);
reg [2055:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1027:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
fsm fsm_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024])); 
fsm fsm_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
fsm fsm_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016])); 
fsm fsm_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
fsm fsm_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
fsm fsm_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013])); 
fsm fsm_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
fsm fsm_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
fsm fsm_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
fsm fsm_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
fsm fsm_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
fsm fsm_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
fsm fsm_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
fsm fsm_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991])); 
fsm fsm_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
mux_module mux_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
mux_module mux_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
fsm fsm_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948])); 
fsm fsm_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
fsm fsm_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
fsm fsm_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
fsm fsm_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
fsm fsm_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
fsm fsm_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935])); 
mux_module mux_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
fsm fsm_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921])); 
fsm fsm_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
fsm fsm_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
fsm fsm_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
fsm fsm_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
mux_module mux_module_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
fsm fsm_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
fsm fsm_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
mux_module mux_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
fsm fsm_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
fsm fsm_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
mux_module mux_module_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
fsm fsm_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
fsm fsm_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
fsm fsm_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
mux_module mux_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
mux_module mux_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
fsm fsm_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
fsm fsm_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865])); 
fsm fsm_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
fsm fsm_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
fsm fsm_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
mux_module mux_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
fsm fsm_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
mux_module mux_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
fsm fsm_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
fsm fsm_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
fsm fsm_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
fsm fsm_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
mux_module mux_module_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
mux_module mux_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
fsm fsm_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
fsm fsm_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
fsm fsm_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
fsm fsm_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
fsm fsm_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
fsm fsm_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
fsm fsm_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
mux_module mux_module_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
mux_module mux_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
mux_module mux_module_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
fsm fsm_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
fsm fsm_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
fsm fsm_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
fsm fsm_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
fsm fsm_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
fsm fsm_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
fsm fsm_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
fsm fsm_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
fsm fsm_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
fsm fsm_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
fsm fsm_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
fsm fsm_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
fsm fsm_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
fsm fsm_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
fsm fsm_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
fsm fsm_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
mux_module mux_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
mux_module mux_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
fsm fsm_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
fsm fsm_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
fsm fsm_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
mux_module mux_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704])); 
fsm fsm_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
fsm fsm_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
fsm fsm_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
fsm fsm_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
mux_module mux_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
fsm fsm_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
mux_module mux_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
fsm fsm_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
mux_module mux_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
fsm fsm_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
mux_module mux_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
fsm fsm_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
mux_module mux_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
fsm fsm_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
fsm fsm_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
mux_module mux_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
fsm fsm_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650])); 
fsm fsm_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
mux_module mux_module_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
fsm fsm_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
fsm fsm_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
fsm fsm_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
mux_module mux_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
mux_module mux_module_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620])); 
fsm fsm_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
fsm fsm_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
mux_module mux_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
mux_module mux_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
fsm fsm_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
mux_module mux_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602])); 
mux_module mux_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600])); 
mux_module mux_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
fsm fsm_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
fsm fsm_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
fsm fsm_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
mux_module mux_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
fsm fsm_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
fsm fsm_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548])); 
fsm fsm_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
mux_module mux_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
fsm fsm_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537])); 
mux_module mux_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
mux_module mux_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
fsm fsm_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
fsm fsm_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
mux_module mux_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513])); 
mux_module mux_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
fsm fsm_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
mux_module mux_module_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
fsm fsm_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
fsm fsm_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
fsm fsm_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
fsm fsm_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
fsm fsm_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
fsm fsm_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
fsm fsm_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
fsm fsm_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
fsm fsm_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
mux_module mux_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
fsm fsm_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
fsm fsm_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
mux_module mux_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
fsm fsm_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
mux_module mux_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
fsm fsm_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
fsm fsm_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
fsm fsm_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
mux_module mux_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
fsm fsm_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
fsm fsm_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
fsm fsm_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
fsm fsm_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
fsm fsm_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
mux_module mux_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
mux_module mux_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
mux_module mux_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
fsm fsm_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
fsm fsm_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
mux_module mux_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
mux_module mux_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
mux_module mux_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
fsm fsm_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
fsm fsm_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
fsm fsm_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
mux_module mux_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
fsm fsm_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
mux_module mux_module_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
fsm fsm_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
fsm fsm_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354])); 
mux_module mux_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
fsm fsm_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
fsm fsm_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
fsm fsm_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
fsm fsm_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
fsm fsm_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
mux_module mux_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
fsm fsm_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338])); 
mux_module mux_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335])); 
fsm fsm_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
fsm fsm_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
fsm fsm_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
fsm fsm_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
fsm fsm_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
mux_module mux_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
mux_module mux_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
fsm fsm_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
fsm fsm_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
fsm fsm_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
fsm fsm_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
fsm fsm_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
fsm fsm_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299])); 
mux_module mux_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
fsm fsm_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
mux_module mux_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
fsm fsm_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
fsm fsm_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
mux_module mux_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
fsm fsm_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
fsm fsm_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
mux_module mux_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
mux_module mux_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
fsm fsm_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
fsm fsm_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
fsm fsm_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
mux_module mux_module_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
fsm fsm_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
mux_module mux_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
fsm fsm_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
mux_module mux_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
mux_module mux_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
mux_module mux_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
fsm fsm_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236])); 
fsm fsm_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
fsm fsm_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
fsm fsm_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
fsm fsm_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
mux_module mux_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
mux_module mux_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
mux_module mux_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221])); 
fsm fsm_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
mux_module mux_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
mux_module mux_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
fsm fsm_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
mux_module mux_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
fsm fsm_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
mux_module mux_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
mux_module mux_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
mux_module mux_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
fsm fsm_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
mux_module mux_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
mux_module mux_module_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
fsm fsm_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
fsm fsm_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
fsm fsm_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
fsm fsm_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
fsm fsm_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
mux_module mux_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
mux_module mux_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
mux_module mux_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
mux_module mux_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
fsm fsm_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
mux_module mux_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
mux_module mux_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
fsm fsm_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
fsm fsm_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
fsm fsm_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
fsm fsm_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
fsm fsm_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
mux_module mux_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
fsm fsm_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
fsm fsm_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
mux_module mux_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
fsm fsm_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
mux_module mux_module_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
mux_module mux_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
fsm fsm_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
mux_module mux_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
mux_module mux_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
mux_module mux_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
mux_module mux_module_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112])); 
fsm fsm_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
mux_module mux_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
fsm fsm_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
mux_module mux_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101])); 
mux_module mux_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
mux_module mux_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
mux_module mux_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82])); 
fsm fsm_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
fsm fsm_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80])); 
mux_module mux_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
mux_module mux_module_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
fsm fsm_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73])); 
fsm fsm_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
mux_module mux_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
fsm fsm_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
mux_module mux_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
fsm fsm_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
fsm fsm_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
fsm fsm_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
mux_module mux_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
mux_module mux_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
fsm fsm_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
mux_module mux_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
mux_module mux_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
fsm fsm_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
mux_module mux_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
fsm fsm_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
fsm fsm_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
mux_module mux_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
fsm fsm_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
mux_module mux_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
fsm fsm_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
mux_module mux_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
mux_module mux_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
fsm fsm_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
fsm fsm_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
fsm fsm_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
mux_module mux_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
mux_module mux_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
fsm fsm_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
fsm fsm_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
fsm fsm_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
mux_module mux_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
mux_module mux_module_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
fsm fsm_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0])); 
reg [513:0]intermediate_reg_2; 
 
fsm fsm_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513])); 
mux_module mux_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510])); 
fsm fsm_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504])); 
fsm fsm_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503])); 
fsm fsm_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502])); 
fsm fsm_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501])); 
fsm fsm_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500])); 
fsm fsm_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499])); 
mux_module mux_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496])); 
fsm fsm_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495])); 
fsm fsm_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494])); 
mux_module mux_module_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491])); 
mux_module mux_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488])); 
mux_module mux_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485])); 
fsm fsm_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484])); 
mux_module mux_module_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
mux_module mux_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477])); 
mux_module mux_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474])); 
mux_module mux_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471])); 
fsm fsm_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470])); 
mux_module mux_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468])); 
fsm fsm_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467])); 
fsm fsm_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466])); 
mux_module mux_module_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464])); 
mux_module mux_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459])); 
fsm fsm_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458])); 
mux_module mux_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456])); 
mux_module mux_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451])); 
mux_module mux_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446])); 
mux_module mux_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443])); 
mux_module mux_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441])); 
mux_module mux_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439])); 
mux_module mux_module_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435])); 
fsm fsm_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434])); 
fsm fsm_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433])); 
fsm fsm_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430])); 
fsm fsm_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429])); 
mux_module mux_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427])); 
mux_module mux_module_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425])); 
fsm fsm_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424])); 
mux_module mux_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420])); 
mux_module mux_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418])); 
mux_module mux_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415])); 
fsm fsm_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414])); 
mux_module mux_module_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412])); 
mux_module mux_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410])); 
mux_module mux_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408])); 
fsm fsm_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407])); 
mux_module mux_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404])); 
mux_module mux_module_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400])); 
mux_module mux_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398])); 
fsm fsm_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397])); 
fsm fsm_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396])); 
mux_module mux_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392])); 
mux_module mux_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387])); 
fsm fsm_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386])); 
fsm fsm_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385])); 
fsm fsm_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384])); 
fsm fsm_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383])); 
mux_module mux_module_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378])); 
fsm fsm_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377])); 
mux_module mux_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375])); 
fsm fsm_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374])); 
fsm fsm_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373])); 
mux_module mux_module_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371])); 
fsm fsm_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
fsm fsm_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369])); 
mux_module mux_module_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367])); 
mux_module mux_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362])); 
fsm fsm_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361])); 
fsm fsm_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360])); 
fsm fsm_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
fsm fsm_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
mux_module mux_module_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356])); 
mux_module mux_module_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354])); 
fsm fsm_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353])); 
mux_module mux_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349])); 
fsm fsm_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348])); 
fsm fsm_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
mux_module mux_module_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
fsm fsm_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343])); 
mux_module mux_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339])); 
fsm fsm_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338])); 
mux_module mux_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
mux_module mux_module_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333])); 
fsm fsm_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332])); 
mux_module mux_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
fsm fsm_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
fsm fsm_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328])); 
fsm fsm_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
mux_module mux_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324])); 
mux_module mux_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322])); 
mux_module mux_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
fsm fsm_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319])); 
mux_module mux_module_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317])); 
mux_module mux_module_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314])); 
fsm fsm_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313])); 
mux_module mux_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311])); 
mux_module mux_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306])); 
mux_module mux_module_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
fsm fsm_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302])); 
fsm fsm_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
fsm fsm_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300])); 
fsm fsm_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299])); 
mux_module mux_module_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297])); 
fsm fsm_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
mux_module mux_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294])); 
fsm fsm_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
mux_module mux_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291])); 
mux_module mux_module_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288])); 
fsm fsm_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287])); 
mux_module mux_module_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
fsm fsm_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284])); 
fsm fsm_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
mux_module mux_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280])); 
mux_module mux_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277])); 
mux_module mux_module_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275])); 
fsm fsm_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
mux_module mux_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269])); 
fsm fsm_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268])); 
mux_module mux_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266])); 
fsm fsm_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
mux_module mux_module_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263])); 
fsm fsm_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
mux_module mux_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259])); 
mux_module mux_module_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257])); 
fsm fsm_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
fsm fsm_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255])); 
mux_module mux_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253])); 
fsm fsm_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252])); 
fsm fsm_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
mux_module mux_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
mux_module mux_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247])); 
fsm fsm_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246])); 
mux_module mux_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
fsm fsm_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240])); 
mux_module mux_module_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
mux_module mux_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234])); 
fsm fsm_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233])); 
mux_module mux_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231])); 
fsm fsm_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230])); 
mux_module mux_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
fsm fsm_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227])); 
mux_module mux_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
mux_module mux_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223])); 
fsm fsm_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
mux_module mux_module_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220])); 
mux_module mux_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
mux_module mux_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
fsm fsm_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
fsm fsm_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
fsm fsm_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
mux_module mux_module_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208])); 
fsm fsm_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
fsm fsm_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
mux_module mux_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204])); 
mux_module mux_module_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201])); 
mux_module mux_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197])); 
fsm fsm_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
mux_module mux_module_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190])); 
mux_module mux_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
mux_module mux_module_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
mux_module mux_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180])); 
mux_module mux_module_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
mux_module mux_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175])); 
mux_module mux_module_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
fsm fsm_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
mux_module mux_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168])); 
mux_module mux_module_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
fsm fsm_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164])); 
fsm fsm_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
fsm fsm_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162])); 
mux_module mux_module_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160])); 
mux_module mux_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158])); 
mux_module mux_module_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155])); 
fsm fsm_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154])); 
fsm fsm_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153])); 
mux_module mux_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
mux_module mux_module_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147])); 
mux_module mux_module_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144])); 
mux_module mux_module_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142])); 
fsm fsm_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141])); 
mux_module mux_module_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139])); 
fsm fsm_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138])); 
mux_module mux_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
mux_module mux_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132])); 
fsm fsm_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131])); 
mux_module mux_module_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
fsm fsm_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
mux_module mux_module_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
mux_module mux_module_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120])); 
mux_module mux_module_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
mux_module mux_module_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
fsm fsm_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
mux_module mux_module_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107])); 
fsm fsm_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
mux_module mux_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104])); 
mux_module mux_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101])); 
mux_module mux_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98])); 
fsm fsm_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
mux_module mux_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94])); 
fsm fsm_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
mux_module mux_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88])); 
mux_module mux_module_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
fsm fsm_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
fsm fsm_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
mux_module mux_module_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82])); 
mux_module mux_module_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77])); 
fsm fsm_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76])); 
mux_module mux_module_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74])); 
mux_module mux_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71])); 
fsm fsm_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
mux_module mux_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66])); 
fsm fsm_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65])); 
mux_module mux_module_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
fsm fsm_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60])); 
mux_module mux_module_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
fsm fsm_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57])); 
fsm fsm_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56])); 
mux_module mux_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
fsm fsm_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
mux_module mux_module_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
mux_module mux_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48])); 
mux_module mux_module_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46])); 
mux_module mux_module_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44])); 
fsm fsm_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
mux_module mux_module_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
mux_module mux_module_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36])); 
fsm fsm_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35])); 
mux_module mux_module_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32])); 
fsm fsm_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
mux_module mux_module_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
mux_module mux_module_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26])); 
mux_module mux_module_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24])); 
mux_module mux_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21])); 
fsm fsm_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20])); 
fsm fsm_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
mux_module mux_module_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17])); 
fsm fsm_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16])); 
mux_module mux_module_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10])); 
mux_module mux_module_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
mux_module mux_module_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
fsm fsm_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0])); 
reg [256:0]intermediate_reg_3; 
 
fsm fsm_inst_3_0(.clk(clk),.reset(reset),.i1(intermediate_reg_2[513]),.i2(intermediate_reg_2[512]),.o(intermediate_reg_3[256])); 
mux_module mux_module_inst_3_1(.clk(clk),.reset(reset),.i1(intermediate_reg_2[511]),.i2(intermediate_reg_2[510]),.o(intermediate_reg_3[255]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_2(.clk(clk),.reset(reset),.i1(intermediate_reg_2[509]),.i2(intermediate_reg_2[508]),.o(intermediate_reg_3[254]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_3(.clk(clk),.reset(reset),.i1(intermediate_reg_2[507]),.i2(intermediate_reg_2[506]),.o(intermediate_reg_3[253])); 
mux_module mux_module_inst_3_4(.clk(clk),.reset(reset),.i1(intermediate_reg_2[505]),.i2(intermediate_reg_2[504]),.o(intermediate_reg_3[252]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_5(.clk(clk),.reset(reset),.i1(intermediate_reg_2[503]),.i2(intermediate_reg_2[502]),.o(intermediate_reg_3[251])); 
mux_module mux_module_inst_3_6(.clk(clk),.reset(reset),.i1(intermediate_reg_2[501]),.i2(intermediate_reg_2[500]),.o(intermediate_reg_3[250]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_7(.clk(clk),.reset(reset),.i1(intermediate_reg_2[499]),.i2(intermediate_reg_2[498]),.o(intermediate_reg_3[249])); 
fsm fsm_inst_3_8(.clk(clk),.reset(reset),.i1(intermediate_reg_2[497]),.i2(intermediate_reg_2[496]),.o(intermediate_reg_3[248])); 
fsm fsm_inst_3_9(.clk(clk),.reset(reset),.i1(intermediate_reg_2[495]),.i2(intermediate_reg_2[494]),.o(intermediate_reg_3[247])); 
mux_module mux_module_inst_3_10(.clk(clk),.reset(reset),.i1(intermediate_reg_2[493]),.i2(intermediate_reg_2[492]),.o(intermediate_reg_3[246]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_11(.clk(clk),.reset(reset),.i1(intermediate_reg_2[491]),.i2(intermediate_reg_2[490]),.o(intermediate_reg_3[245]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_12(.clk(clk),.reset(reset),.i1(intermediate_reg_2[489]),.i2(intermediate_reg_2[488]),.o(intermediate_reg_3[244])); 
mux_module mux_module_inst_3_13(.clk(clk),.reset(reset),.i1(intermediate_reg_2[487]),.i2(intermediate_reg_2[486]),.o(intermediate_reg_3[243]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_14(.clk(clk),.reset(reset),.i1(intermediate_reg_2[485]),.i2(intermediate_reg_2[484]),.o(intermediate_reg_3[242]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_15(.clk(clk),.reset(reset),.i1(intermediate_reg_2[483]),.i2(intermediate_reg_2[482]),.o(intermediate_reg_3[241])); 
fsm fsm_inst_3_16(.clk(clk),.reset(reset),.i1(intermediate_reg_2[481]),.i2(intermediate_reg_2[480]),.o(intermediate_reg_3[240])); 
fsm fsm_inst_3_17(.clk(clk),.reset(reset),.i1(intermediate_reg_2[479]),.i2(intermediate_reg_2[478]),.o(intermediate_reg_3[239])); 
fsm fsm_inst_3_18(.clk(clk),.reset(reset),.i1(intermediate_reg_2[477]),.i2(intermediate_reg_2[476]),.o(intermediate_reg_3[238])); 
fsm fsm_inst_3_19(.clk(clk),.reset(reset),.i1(intermediate_reg_2[475]),.i2(intermediate_reg_2[474]),.o(intermediate_reg_3[237])); 
mux_module mux_module_inst_3_20(.clk(clk),.reset(reset),.i1(intermediate_reg_2[473]),.i2(intermediate_reg_2[472]),.o(intermediate_reg_3[236]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_21(.clk(clk),.reset(reset),.i1(intermediate_reg_2[471]),.i2(intermediate_reg_2[470]),.o(intermediate_reg_3[235]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_22(.clk(clk),.reset(reset),.i1(intermediate_reg_2[469]),.i2(intermediate_reg_2[468]),.o(intermediate_reg_3[234]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_23(.clk(clk),.reset(reset),.i1(intermediate_reg_2[467]),.i2(intermediate_reg_2[466]),.o(intermediate_reg_3[233]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_24(.clk(clk),.reset(reset),.i1(intermediate_reg_2[465]),.i2(intermediate_reg_2[464]),.o(intermediate_reg_3[232]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_25(.clk(clk),.reset(reset),.i1(intermediate_reg_2[463]),.i2(intermediate_reg_2[462]),.o(intermediate_reg_3[231]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_26(.clk(clk),.reset(reset),.i1(intermediate_reg_2[461]),.i2(intermediate_reg_2[460]),.o(intermediate_reg_3[230])); 
fsm fsm_inst_3_27(.clk(clk),.reset(reset),.i1(intermediate_reg_2[459]),.i2(intermediate_reg_2[458]),.o(intermediate_reg_3[229])); 
fsm fsm_inst_3_28(.clk(clk),.reset(reset),.i1(intermediate_reg_2[457]),.i2(intermediate_reg_2[456]),.o(intermediate_reg_3[228])); 
fsm fsm_inst_3_29(.clk(clk),.reset(reset),.i1(intermediate_reg_2[455]),.i2(intermediate_reg_2[454]),.o(intermediate_reg_3[227])); 
mux_module mux_module_inst_3_30(.clk(clk),.reset(reset),.i1(intermediate_reg_2[453]),.i2(intermediate_reg_2[452]),.o(intermediate_reg_3[226]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_31(.clk(clk),.reset(reset),.i1(intermediate_reg_2[451]),.i2(intermediate_reg_2[450]),.o(intermediate_reg_3[225]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_32(.clk(clk),.reset(reset),.i1(intermediate_reg_2[449]),.i2(intermediate_reg_2[448]),.o(intermediate_reg_3[224]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_33(.clk(clk),.reset(reset),.i1(intermediate_reg_2[447]),.i2(intermediate_reg_2[446]),.o(intermediate_reg_3[223])); 
fsm fsm_inst_3_34(.clk(clk),.reset(reset),.i1(intermediate_reg_2[445]),.i2(intermediate_reg_2[444]),.o(intermediate_reg_3[222])); 
mux_module mux_module_inst_3_35(.clk(clk),.reset(reset),.i1(intermediate_reg_2[443]),.i2(intermediate_reg_2[442]),.o(intermediate_reg_3[221]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_36(.clk(clk),.reset(reset),.i1(intermediate_reg_2[441]),.i2(intermediate_reg_2[440]),.o(intermediate_reg_3[220]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_37(.clk(clk),.reset(reset),.i1(intermediate_reg_2[439]),.i2(intermediate_reg_2[438]),.o(intermediate_reg_3[219])); 
mux_module mux_module_inst_3_38(.clk(clk),.reset(reset),.i1(intermediate_reg_2[437]),.i2(intermediate_reg_2[436]),.o(intermediate_reg_3[218]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_39(.clk(clk),.reset(reset),.i1(intermediate_reg_2[435]),.i2(intermediate_reg_2[434]),.o(intermediate_reg_3[217])); 
fsm fsm_inst_3_40(.clk(clk),.reset(reset),.i1(intermediate_reg_2[433]),.i2(intermediate_reg_2[432]),.o(intermediate_reg_3[216])); 
fsm fsm_inst_3_41(.clk(clk),.reset(reset),.i1(intermediate_reg_2[431]),.i2(intermediate_reg_2[430]),.o(intermediate_reg_3[215])); 
fsm fsm_inst_3_42(.clk(clk),.reset(reset),.i1(intermediate_reg_2[429]),.i2(intermediate_reg_2[428]),.o(intermediate_reg_3[214])); 
mux_module mux_module_inst_3_43(.clk(clk),.reset(reset),.i1(intermediate_reg_2[427]),.i2(intermediate_reg_2[426]),.o(intermediate_reg_3[213]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_44(.clk(clk),.reset(reset),.i1(intermediate_reg_2[425]),.i2(intermediate_reg_2[424]),.o(intermediate_reg_3[212]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_45(.clk(clk),.reset(reset),.i1(intermediate_reg_2[423]),.i2(intermediate_reg_2[422]),.o(intermediate_reg_3[211]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_46(.clk(clk),.reset(reset),.i1(intermediate_reg_2[421]),.i2(intermediate_reg_2[420]),.o(intermediate_reg_3[210])); 
mux_module mux_module_inst_3_47(.clk(clk),.reset(reset),.i1(intermediate_reg_2[419]),.i2(intermediate_reg_2[418]),.o(intermediate_reg_3[209]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_48(.clk(clk),.reset(reset),.i1(intermediate_reg_2[417]),.i2(intermediate_reg_2[416]),.o(intermediate_reg_3[208]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_49(.clk(clk),.reset(reset),.i1(intermediate_reg_2[415]),.i2(intermediate_reg_2[414]),.o(intermediate_reg_3[207])); 
fsm fsm_inst_3_50(.clk(clk),.reset(reset),.i1(intermediate_reg_2[413]),.i2(intermediate_reg_2[412]),.o(intermediate_reg_3[206])); 
mux_module mux_module_inst_3_51(.clk(clk),.reset(reset),.i1(intermediate_reg_2[411]),.i2(intermediate_reg_2[410]),.o(intermediate_reg_3[205]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_52(.clk(clk),.reset(reset),.i1(intermediate_reg_2[409]),.i2(intermediate_reg_2[408]),.o(intermediate_reg_3[204]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_53(.clk(clk),.reset(reset),.i1(intermediate_reg_2[407]),.i2(intermediate_reg_2[406]),.o(intermediate_reg_3[203]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_54(.clk(clk),.reset(reset),.i1(intermediate_reg_2[405]),.i2(intermediate_reg_2[404]),.o(intermediate_reg_3[202])); 
fsm fsm_inst_3_55(.clk(clk),.reset(reset),.i1(intermediate_reg_2[403]),.i2(intermediate_reg_2[402]),.o(intermediate_reg_3[201])); 
mux_module mux_module_inst_3_56(.clk(clk),.reset(reset),.i1(intermediate_reg_2[401]),.i2(intermediate_reg_2[400]),.o(intermediate_reg_3[200]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_57(.clk(clk),.reset(reset),.i1(intermediate_reg_2[399]),.i2(intermediate_reg_2[398]),.o(intermediate_reg_3[199])); 
mux_module mux_module_inst_3_58(.clk(clk),.reset(reset),.i1(intermediate_reg_2[397]),.i2(intermediate_reg_2[396]),.o(intermediate_reg_3[198]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_59(.clk(clk),.reset(reset),.i1(intermediate_reg_2[395]),.i2(intermediate_reg_2[394]),.o(intermediate_reg_3[197]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_60(.clk(clk),.reset(reset),.i1(intermediate_reg_2[393]),.i2(intermediate_reg_2[392]),.o(intermediate_reg_3[196])); 
mux_module mux_module_inst_3_61(.clk(clk),.reset(reset),.i1(intermediate_reg_2[391]),.i2(intermediate_reg_2[390]),.o(intermediate_reg_3[195]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_62(.clk(clk),.reset(reset),.i1(intermediate_reg_2[389]),.i2(intermediate_reg_2[388]),.o(intermediate_reg_3[194])); 
fsm fsm_inst_3_63(.clk(clk),.reset(reset),.i1(intermediate_reg_2[387]),.i2(intermediate_reg_2[386]),.o(intermediate_reg_3[193])); 
fsm fsm_inst_3_64(.clk(clk),.reset(reset),.i1(intermediate_reg_2[385]),.i2(intermediate_reg_2[384]),.o(intermediate_reg_3[192])); 
fsm fsm_inst_3_65(.clk(clk),.reset(reset),.i1(intermediate_reg_2[383]),.i2(intermediate_reg_2[382]),.o(intermediate_reg_3[191])); 
fsm fsm_inst_3_66(.clk(clk),.reset(reset),.i1(intermediate_reg_2[381]),.i2(intermediate_reg_2[380]),.o(intermediate_reg_3[190])); 
mux_module mux_module_inst_3_67(.clk(clk),.reset(reset),.i1(intermediate_reg_2[379]),.i2(intermediate_reg_2[378]),.o(intermediate_reg_3[189]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_68(.clk(clk),.reset(reset),.i1(intermediate_reg_2[377]),.i2(intermediate_reg_2[376]),.o(intermediate_reg_3[188])); 
mux_module mux_module_inst_3_69(.clk(clk),.reset(reset),.i1(intermediate_reg_2[375]),.i2(intermediate_reg_2[374]),.o(intermediate_reg_3[187]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_70(.clk(clk),.reset(reset),.i1(intermediate_reg_2[373]),.i2(intermediate_reg_2[372]),.o(intermediate_reg_3[186])); 
mux_module mux_module_inst_3_71(.clk(clk),.reset(reset),.i1(intermediate_reg_2[371]),.i2(intermediate_reg_2[370]),.o(intermediate_reg_3[185]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_72(.clk(clk),.reset(reset),.i1(intermediate_reg_2[369]),.i2(intermediate_reg_2[368]),.o(intermediate_reg_3[184])); 
fsm fsm_inst_3_73(.clk(clk),.reset(reset),.i1(intermediate_reg_2[367]),.i2(intermediate_reg_2[366]),.o(intermediate_reg_3[183])); 
fsm fsm_inst_3_74(.clk(clk),.reset(reset),.i1(intermediate_reg_2[365]),.i2(intermediate_reg_2[364]),.o(intermediate_reg_3[182])); 
fsm fsm_inst_3_75(.clk(clk),.reset(reset),.i1(intermediate_reg_2[363]),.i2(intermediate_reg_2[362]),.o(intermediate_reg_3[181])); 
mux_module mux_module_inst_3_76(.clk(clk),.reset(reset),.i1(intermediate_reg_2[361]),.i2(intermediate_reg_2[360]),.o(intermediate_reg_3[180]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_77(.clk(clk),.reset(reset),.i1(intermediate_reg_2[359]),.i2(intermediate_reg_2[358]),.o(intermediate_reg_3[179]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_78(.clk(clk),.reset(reset),.i1(intermediate_reg_2[357]),.i2(intermediate_reg_2[356]),.o(intermediate_reg_3[178])); 
fsm fsm_inst_3_79(.clk(clk),.reset(reset),.i1(intermediate_reg_2[355]),.i2(intermediate_reg_2[354]),.o(intermediate_reg_3[177])); 
fsm fsm_inst_3_80(.clk(clk),.reset(reset),.i1(intermediate_reg_2[353]),.i2(intermediate_reg_2[352]),.o(intermediate_reg_3[176])); 
fsm fsm_inst_3_81(.clk(clk),.reset(reset),.i1(intermediate_reg_2[351]),.i2(intermediate_reg_2[350]),.o(intermediate_reg_3[175])); 
mux_module mux_module_inst_3_82(.clk(clk),.reset(reset),.i1(intermediate_reg_2[349]),.i2(intermediate_reg_2[348]),.o(intermediate_reg_3[174]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_83(.clk(clk),.reset(reset),.i1(intermediate_reg_2[347]),.i2(intermediate_reg_2[346]),.o(intermediate_reg_3[173]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_84(.clk(clk),.reset(reset),.i1(intermediate_reg_2[345]),.i2(intermediate_reg_2[344]),.o(intermediate_reg_3[172])); 
fsm fsm_inst_3_85(.clk(clk),.reset(reset),.i1(intermediate_reg_2[343]),.i2(intermediate_reg_2[342]),.o(intermediate_reg_3[171])); 
mux_module mux_module_inst_3_86(.clk(clk),.reset(reset),.i1(intermediate_reg_2[341]),.i2(intermediate_reg_2[340]),.o(intermediate_reg_3[170]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_87(.clk(clk),.reset(reset),.i1(intermediate_reg_2[339]),.i2(intermediate_reg_2[338]),.o(intermediate_reg_3[169]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_88(.clk(clk),.reset(reset),.i1(intermediate_reg_2[337]),.i2(intermediate_reg_2[336]),.o(intermediate_reg_3[168]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_89(.clk(clk),.reset(reset),.i1(intermediate_reg_2[335]),.i2(intermediate_reg_2[334]),.o(intermediate_reg_3[167]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_90(.clk(clk),.reset(reset),.i1(intermediate_reg_2[333]),.i2(intermediate_reg_2[332]),.o(intermediate_reg_3[166]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_91(.clk(clk),.reset(reset),.i1(intermediate_reg_2[331]),.i2(intermediate_reg_2[330]),.o(intermediate_reg_3[165]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_92(.clk(clk),.reset(reset),.i1(intermediate_reg_2[329]),.i2(intermediate_reg_2[328]),.o(intermediate_reg_3[164]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_93(.clk(clk),.reset(reset),.i1(intermediate_reg_2[327]),.i2(intermediate_reg_2[326]),.o(intermediate_reg_3[163])); 
mux_module mux_module_inst_3_94(.clk(clk),.reset(reset),.i1(intermediate_reg_2[325]),.i2(intermediate_reg_2[324]),.o(intermediate_reg_3[162]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_95(.clk(clk),.reset(reset),.i1(intermediate_reg_2[323]),.i2(intermediate_reg_2[322]),.o(intermediate_reg_3[161]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_96(.clk(clk),.reset(reset),.i1(intermediate_reg_2[321]),.i2(intermediate_reg_2[320]),.o(intermediate_reg_3[160]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_97(.clk(clk),.reset(reset),.i1(intermediate_reg_2[319]),.i2(intermediate_reg_2[318]),.o(intermediate_reg_3[159]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_98(.clk(clk),.reset(reset),.i1(intermediate_reg_2[317]),.i2(intermediate_reg_2[316]),.o(intermediate_reg_3[158]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_99(.clk(clk),.reset(reset),.i1(intermediate_reg_2[315]),.i2(intermediate_reg_2[314]),.o(intermediate_reg_3[157])); 
mux_module mux_module_inst_3_100(.clk(clk),.reset(reset),.i1(intermediate_reg_2[313]),.i2(intermediate_reg_2[312]),.o(intermediate_reg_3[156]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_101(.clk(clk),.reset(reset),.i1(intermediate_reg_2[311]),.i2(intermediate_reg_2[310]),.o(intermediate_reg_3[155])); 
mux_module mux_module_inst_3_102(.clk(clk),.reset(reset),.i1(intermediate_reg_2[309]),.i2(intermediate_reg_2[308]),.o(intermediate_reg_3[154]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_103(.clk(clk),.reset(reset),.i1(intermediate_reg_2[307]),.i2(intermediate_reg_2[306]),.o(intermediate_reg_3[153]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_104(.clk(clk),.reset(reset),.i1(intermediate_reg_2[305]),.i2(intermediate_reg_2[304]),.o(intermediate_reg_3[152]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_105(.clk(clk),.reset(reset),.i1(intermediate_reg_2[303]),.i2(intermediate_reg_2[302]),.o(intermediate_reg_3[151])); 
fsm fsm_inst_3_106(.clk(clk),.reset(reset),.i1(intermediate_reg_2[301]),.i2(intermediate_reg_2[300]),.o(intermediate_reg_3[150])); 
mux_module mux_module_inst_3_107(.clk(clk),.reset(reset),.i1(intermediate_reg_2[299]),.i2(intermediate_reg_2[298]),.o(intermediate_reg_3[149]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_108(.clk(clk),.reset(reset),.i1(intermediate_reg_2[297]),.i2(intermediate_reg_2[296]),.o(intermediate_reg_3[148]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_109(.clk(clk),.reset(reset),.i1(intermediate_reg_2[295]),.i2(intermediate_reg_2[294]),.o(intermediate_reg_3[147])); 
mux_module mux_module_inst_3_110(.clk(clk),.reset(reset),.i1(intermediate_reg_2[293]),.i2(intermediate_reg_2[292]),.o(intermediate_reg_3[146]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_111(.clk(clk),.reset(reset),.i1(intermediate_reg_2[291]),.i2(intermediate_reg_2[290]),.o(intermediate_reg_3[145]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_112(.clk(clk),.reset(reset),.i1(intermediate_reg_2[289]),.i2(intermediate_reg_2[288]),.o(intermediate_reg_3[144])); 
fsm fsm_inst_3_113(.clk(clk),.reset(reset),.i1(intermediate_reg_2[287]),.i2(intermediate_reg_2[286]),.o(intermediate_reg_3[143])); 
fsm fsm_inst_3_114(.clk(clk),.reset(reset),.i1(intermediate_reg_2[285]),.i2(intermediate_reg_2[284]),.o(intermediate_reg_3[142])); 
mux_module mux_module_inst_3_115(.clk(clk),.reset(reset),.i1(intermediate_reg_2[283]),.i2(intermediate_reg_2[282]),.o(intermediate_reg_3[141]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_116(.clk(clk),.reset(reset),.i1(intermediate_reg_2[281]),.i2(intermediate_reg_2[280]),.o(intermediate_reg_3[140]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_117(.clk(clk),.reset(reset),.i1(intermediate_reg_2[279]),.i2(intermediate_reg_2[278]),.o(intermediate_reg_3[139]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_118(.clk(clk),.reset(reset),.i1(intermediate_reg_2[277]),.i2(intermediate_reg_2[276]),.o(intermediate_reg_3[138]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_119(.clk(clk),.reset(reset),.i1(intermediate_reg_2[275]),.i2(intermediate_reg_2[274]),.o(intermediate_reg_3[137]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_120(.clk(clk),.reset(reset),.i1(intermediate_reg_2[273]),.i2(intermediate_reg_2[272]),.o(intermediate_reg_3[136])); 
mux_module mux_module_inst_3_121(.clk(clk),.reset(reset),.i1(intermediate_reg_2[271]),.i2(intermediate_reg_2[270]),.o(intermediate_reg_3[135]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_122(.clk(clk),.reset(reset),.i1(intermediate_reg_2[269]),.i2(intermediate_reg_2[268]),.o(intermediate_reg_3[134]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_123(.clk(clk),.reset(reset),.i1(intermediate_reg_2[267]),.i2(intermediate_reg_2[266]),.o(intermediate_reg_3[133]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_124(.clk(clk),.reset(reset),.i1(intermediate_reg_2[265]),.i2(intermediate_reg_2[264]),.o(intermediate_reg_3[132])); 
fsm fsm_inst_3_125(.clk(clk),.reset(reset),.i1(intermediate_reg_2[263]),.i2(intermediate_reg_2[262]),.o(intermediate_reg_3[131])); 
mux_module mux_module_inst_3_126(.clk(clk),.reset(reset),.i1(intermediate_reg_2[261]),.i2(intermediate_reg_2[260]),.o(intermediate_reg_3[130]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_127(.clk(clk),.reset(reset),.i1(intermediate_reg_2[259]),.i2(intermediate_reg_2[258]),.o(intermediate_reg_3[129])); 
mux_module mux_module_inst_3_128(.clk(clk),.reset(reset),.i1(intermediate_reg_2[257]),.i2(intermediate_reg_2[256]),.o(intermediate_reg_3[128]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_129(.clk(clk),.reset(reset),.i1(intermediate_reg_2[255]),.i2(intermediate_reg_2[254]),.o(intermediate_reg_3[127])); 
fsm fsm_inst_3_130(.clk(clk),.reset(reset),.i1(intermediate_reg_2[253]),.i2(intermediate_reg_2[252]),.o(intermediate_reg_3[126])); 
fsm fsm_inst_3_131(.clk(clk),.reset(reset),.i1(intermediate_reg_2[251]),.i2(intermediate_reg_2[250]),.o(intermediate_reg_3[125])); 
fsm fsm_inst_3_132(.clk(clk),.reset(reset),.i1(intermediate_reg_2[249]),.i2(intermediate_reg_2[248]),.o(intermediate_reg_3[124])); 
fsm fsm_inst_3_133(.clk(clk),.reset(reset),.i1(intermediate_reg_2[247]),.i2(intermediate_reg_2[246]),.o(intermediate_reg_3[123])); 
fsm fsm_inst_3_134(.clk(clk),.reset(reset),.i1(intermediate_reg_2[245]),.i2(intermediate_reg_2[244]),.o(intermediate_reg_3[122])); 
fsm fsm_inst_3_135(.clk(clk),.reset(reset),.i1(intermediate_reg_2[243]),.i2(intermediate_reg_2[242]),.o(intermediate_reg_3[121])); 
fsm fsm_inst_3_136(.clk(clk),.reset(reset),.i1(intermediate_reg_2[241]),.i2(intermediate_reg_2[240]),.o(intermediate_reg_3[120])); 
mux_module mux_module_inst_3_137(.clk(clk),.reset(reset),.i1(intermediate_reg_2[239]),.i2(intermediate_reg_2[238]),.o(intermediate_reg_3[119]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_138(.clk(clk),.reset(reset),.i1(intermediate_reg_2[237]),.i2(intermediate_reg_2[236]),.o(intermediate_reg_3[118])); 
fsm fsm_inst_3_139(.clk(clk),.reset(reset),.i1(intermediate_reg_2[235]),.i2(intermediate_reg_2[234]),.o(intermediate_reg_3[117])); 
mux_module mux_module_inst_3_140(.clk(clk),.reset(reset),.i1(intermediate_reg_2[233]),.i2(intermediate_reg_2[232]),.o(intermediate_reg_3[116]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_141(.clk(clk),.reset(reset),.i1(intermediate_reg_2[231]),.i2(intermediate_reg_2[230]),.o(intermediate_reg_3[115])); 
mux_module mux_module_inst_3_142(.clk(clk),.reset(reset),.i1(intermediate_reg_2[229]),.i2(intermediate_reg_2[228]),.o(intermediate_reg_3[114]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_143(.clk(clk),.reset(reset),.i1(intermediate_reg_2[227]),.i2(intermediate_reg_2[226]),.o(intermediate_reg_3[113])); 
mux_module mux_module_inst_3_144(.clk(clk),.reset(reset),.i1(intermediate_reg_2[225]),.i2(intermediate_reg_2[224]),.o(intermediate_reg_3[112]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_145(.clk(clk),.reset(reset),.i1(intermediate_reg_2[223]),.i2(intermediate_reg_2[222]),.o(intermediate_reg_3[111]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_146(.clk(clk),.reset(reset),.i1(intermediate_reg_2[221]),.i2(intermediate_reg_2[220]),.o(intermediate_reg_3[110]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_147(.clk(clk),.reset(reset),.i1(intermediate_reg_2[219]),.i2(intermediate_reg_2[218]),.o(intermediate_reg_3[109]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_148(.clk(clk),.reset(reset),.i1(intermediate_reg_2[217]),.i2(intermediate_reg_2[216]),.o(intermediate_reg_3[108])); 
fsm fsm_inst_3_149(.clk(clk),.reset(reset),.i1(intermediate_reg_2[215]),.i2(intermediate_reg_2[214]),.o(intermediate_reg_3[107])); 
fsm fsm_inst_3_150(.clk(clk),.reset(reset),.i1(intermediate_reg_2[213]),.i2(intermediate_reg_2[212]),.o(intermediate_reg_3[106])); 
mux_module mux_module_inst_3_151(.clk(clk),.reset(reset),.i1(intermediate_reg_2[211]),.i2(intermediate_reg_2[210]),.o(intermediate_reg_3[105]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_152(.clk(clk),.reset(reset),.i1(intermediate_reg_2[209]),.i2(intermediate_reg_2[208]),.o(intermediate_reg_3[104]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_153(.clk(clk),.reset(reset),.i1(intermediate_reg_2[207]),.i2(intermediate_reg_2[206]),.o(intermediate_reg_3[103]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_154(.clk(clk),.reset(reset),.i1(intermediate_reg_2[205]),.i2(intermediate_reg_2[204]),.o(intermediate_reg_3[102]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_155(.clk(clk),.reset(reset),.i1(intermediate_reg_2[203]),.i2(intermediate_reg_2[202]),.o(intermediate_reg_3[101]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_156(.clk(clk),.reset(reset),.i1(intermediate_reg_2[201]),.i2(intermediate_reg_2[200]),.o(intermediate_reg_3[100])); 
mux_module mux_module_inst_3_157(.clk(clk),.reset(reset),.i1(intermediate_reg_2[199]),.i2(intermediate_reg_2[198]),.o(intermediate_reg_3[99]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_158(.clk(clk),.reset(reset),.i1(intermediate_reg_2[197]),.i2(intermediate_reg_2[196]),.o(intermediate_reg_3[98]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_159(.clk(clk),.reset(reset),.i1(intermediate_reg_2[195]),.i2(intermediate_reg_2[194]),.o(intermediate_reg_3[97]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_160(.clk(clk),.reset(reset),.i1(intermediate_reg_2[193]),.i2(intermediate_reg_2[192]),.o(intermediate_reg_3[96]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_161(.clk(clk),.reset(reset),.i1(intermediate_reg_2[191]),.i2(intermediate_reg_2[190]),.o(intermediate_reg_3[95])); 
fsm fsm_inst_3_162(.clk(clk),.reset(reset),.i1(intermediate_reg_2[189]),.i2(intermediate_reg_2[188]),.o(intermediate_reg_3[94])); 
fsm fsm_inst_3_163(.clk(clk),.reset(reset),.i1(intermediate_reg_2[187]),.i2(intermediate_reg_2[186]),.o(intermediate_reg_3[93])); 
fsm fsm_inst_3_164(.clk(clk),.reset(reset),.i1(intermediate_reg_2[185]),.i2(intermediate_reg_2[184]),.o(intermediate_reg_3[92])); 
mux_module mux_module_inst_3_165(.clk(clk),.reset(reset),.i1(intermediate_reg_2[183]),.i2(intermediate_reg_2[182]),.o(intermediate_reg_3[91]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_166(.clk(clk),.reset(reset),.i1(intermediate_reg_2[181]),.i2(intermediate_reg_2[180]),.o(intermediate_reg_3[90])); 
mux_module mux_module_inst_3_167(.clk(clk),.reset(reset),.i1(intermediate_reg_2[179]),.i2(intermediate_reg_2[178]),.o(intermediate_reg_3[89]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_168(.clk(clk),.reset(reset),.i1(intermediate_reg_2[177]),.i2(intermediate_reg_2[176]),.o(intermediate_reg_3[88])); 
fsm fsm_inst_3_169(.clk(clk),.reset(reset),.i1(intermediate_reg_2[175]),.i2(intermediate_reg_2[174]),.o(intermediate_reg_3[87])); 
fsm fsm_inst_3_170(.clk(clk),.reset(reset),.i1(intermediate_reg_2[173]),.i2(intermediate_reg_2[172]),.o(intermediate_reg_3[86])); 
fsm fsm_inst_3_171(.clk(clk),.reset(reset),.i1(intermediate_reg_2[171]),.i2(intermediate_reg_2[170]),.o(intermediate_reg_3[85])); 
fsm fsm_inst_3_172(.clk(clk),.reset(reset),.i1(intermediate_reg_2[169]),.i2(intermediate_reg_2[168]),.o(intermediate_reg_3[84])); 
fsm fsm_inst_3_173(.clk(clk),.reset(reset),.i1(intermediate_reg_2[167]),.i2(intermediate_reg_2[166]),.o(intermediate_reg_3[83])); 
fsm fsm_inst_3_174(.clk(clk),.reset(reset),.i1(intermediate_reg_2[165]),.i2(intermediate_reg_2[164]),.o(intermediate_reg_3[82])); 
mux_module mux_module_inst_3_175(.clk(clk),.reset(reset),.i1(intermediate_reg_2[163]),.i2(intermediate_reg_2[162]),.o(intermediate_reg_3[81]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_176(.clk(clk),.reset(reset),.i1(intermediate_reg_2[161]),.i2(intermediate_reg_2[160]),.o(intermediate_reg_3[80])); 
fsm fsm_inst_3_177(.clk(clk),.reset(reset),.i1(intermediate_reg_2[159]),.i2(intermediate_reg_2[158]),.o(intermediate_reg_3[79])); 
fsm fsm_inst_3_178(.clk(clk),.reset(reset),.i1(intermediate_reg_2[157]),.i2(intermediate_reg_2[156]),.o(intermediate_reg_3[78])); 
fsm fsm_inst_3_179(.clk(clk),.reset(reset),.i1(intermediate_reg_2[155]),.i2(intermediate_reg_2[154]),.o(intermediate_reg_3[77])); 
fsm fsm_inst_3_180(.clk(clk),.reset(reset),.i1(intermediate_reg_2[153]),.i2(intermediate_reg_2[152]),.o(intermediate_reg_3[76])); 
mux_module mux_module_inst_3_181(.clk(clk),.reset(reset),.i1(intermediate_reg_2[151]),.i2(intermediate_reg_2[150]),.o(intermediate_reg_3[75]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_182(.clk(clk),.reset(reset),.i1(intermediate_reg_2[149]),.i2(intermediate_reg_2[148]),.o(intermediate_reg_3[74])); 
fsm fsm_inst_3_183(.clk(clk),.reset(reset),.i1(intermediate_reg_2[147]),.i2(intermediate_reg_2[146]),.o(intermediate_reg_3[73])); 
mux_module mux_module_inst_3_184(.clk(clk),.reset(reset),.i1(intermediate_reg_2[145]),.i2(intermediate_reg_2[144]),.o(intermediate_reg_3[72]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_185(.clk(clk),.reset(reset),.i1(intermediate_reg_2[143]),.i2(intermediate_reg_2[142]),.o(intermediate_reg_3[71])); 
mux_module mux_module_inst_3_186(.clk(clk),.reset(reset),.i1(intermediate_reg_2[141]),.i2(intermediate_reg_2[140]),.o(intermediate_reg_3[70]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_187(.clk(clk),.reset(reset),.i1(intermediate_reg_2[139]),.i2(intermediate_reg_2[138]),.o(intermediate_reg_3[69]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_188(.clk(clk),.reset(reset),.i1(intermediate_reg_2[137]),.i2(intermediate_reg_2[136]),.o(intermediate_reg_3[68])); 
mux_module mux_module_inst_3_189(.clk(clk),.reset(reset),.i1(intermediate_reg_2[135]),.i2(intermediate_reg_2[134]),.o(intermediate_reg_3[67]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_190(.clk(clk),.reset(reset),.i1(intermediate_reg_2[133]),.i2(intermediate_reg_2[132]),.o(intermediate_reg_3[66])); 
fsm fsm_inst_3_191(.clk(clk),.reset(reset),.i1(intermediate_reg_2[131]),.i2(intermediate_reg_2[130]),.o(intermediate_reg_3[65])); 
mux_module mux_module_inst_3_192(.clk(clk),.reset(reset),.i1(intermediate_reg_2[129]),.i2(intermediate_reg_2[128]),.o(intermediate_reg_3[64]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_193(.clk(clk),.reset(reset),.i1(intermediate_reg_2[127]),.i2(intermediate_reg_2[126]),.o(intermediate_reg_3[63]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_194(.clk(clk),.reset(reset),.i1(intermediate_reg_2[125]),.i2(intermediate_reg_2[124]),.o(intermediate_reg_3[62]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_195(.clk(clk),.reset(reset),.i1(intermediate_reg_2[123]),.i2(intermediate_reg_2[122]),.o(intermediate_reg_3[61]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_196(.clk(clk),.reset(reset),.i1(intermediate_reg_2[121]),.i2(intermediate_reg_2[120]),.o(intermediate_reg_3[60]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_197(.clk(clk),.reset(reset),.i1(intermediate_reg_2[119]),.i2(intermediate_reg_2[118]),.o(intermediate_reg_3[59])); 
mux_module mux_module_inst_3_198(.clk(clk),.reset(reset),.i1(intermediate_reg_2[117]),.i2(intermediate_reg_2[116]),.o(intermediate_reg_3[58]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_199(.clk(clk),.reset(reset),.i1(intermediate_reg_2[115]),.i2(intermediate_reg_2[114]),.o(intermediate_reg_3[57]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_200(.clk(clk),.reset(reset),.i1(intermediate_reg_2[113]),.i2(intermediate_reg_2[112]),.o(intermediate_reg_3[56]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_201(.clk(clk),.reset(reset),.i1(intermediate_reg_2[111]),.i2(intermediate_reg_2[110]),.o(intermediate_reg_3[55]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_202(.clk(clk),.reset(reset),.i1(intermediate_reg_2[109]),.i2(intermediate_reg_2[108]),.o(intermediate_reg_3[54]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_203(.clk(clk),.reset(reset),.i1(intermediate_reg_2[107]),.i2(intermediate_reg_2[106]),.o(intermediate_reg_3[53])); 
mux_module mux_module_inst_3_204(.clk(clk),.reset(reset),.i1(intermediate_reg_2[105]),.i2(intermediate_reg_2[104]),.o(intermediate_reg_3[52]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_205(.clk(clk),.reset(reset),.i1(intermediate_reg_2[103]),.i2(intermediate_reg_2[102]),.o(intermediate_reg_3[51])); 
fsm fsm_inst_3_206(.clk(clk),.reset(reset),.i1(intermediate_reg_2[101]),.i2(intermediate_reg_2[100]),.o(intermediate_reg_3[50])); 
fsm fsm_inst_3_207(.clk(clk),.reset(reset),.i1(intermediate_reg_2[99]),.i2(intermediate_reg_2[98]),.o(intermediate_reg_3[49])); 
fsm fsm_inst_3_208(.clk(clk),.reset(reset),.i1(intermediate_reg_2[97]),.i2(intermediate_reg_2[96]),.o(intermediate_reg_3[48])); 
mux_module mux_module_inst_3_209(.clk(clk),.reset(reset),.i1(intermediate_reg_2[95]),.i2(intermediate_reg_2[94]),.o(intermediate_reg_3[47]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_210(.clk(clk),.reset(reset),.i1(intermediate_reg_2[93]),.i2(intermediate_reg_2[92]),.o(intermediate_reg_3[46]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_211(.clk(clk),.reset(reset),.i1(intermediate_reg_2[91]),.i2(intermediate_reg_2[90]),.o(intermediate_reg_3[45]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_212(.clk(clk),.reset(reset),.i1(intermediate_reg_2[89]),.i2(intermediate_reg_2[88]),.o(intermediate_reg_3[44])); 
fsm fsm_inst_3_213(.clk(clk),.reset(reset),.i1(intermediate_reg_2[87]),.i2(intermediate_reg_2[86]),.o(intermediate_reg_3[43])); 
fsm fsm_inst_3_214(.clk(clk),.reset(reset),.i1(intermediate_reg_2[85]),.i2(intermediate_reg_2[84]),.o(intermediate_reg_3[42])); 
mux_module mux_module_inst_3_215(.clk(clk),.reset(reset),.i1(intermediate_reg_2[83]),.i2(intermediate_reg_2[82]),.o(intermediate_reg_3[41]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_216(.clk(clk),.reset(reset),.i1(intermediate_reg_2[81]),.i2(intermediate_reg_2[80]),.o(intermediate_reg_3[40]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_217(.clk(clk),.reset(reset),.i1(intermediate_reg_2[79]),.i2(intermediate_reg_2[78]),.o(intermediate_reg_3[39])); 
fsm fsm_inst_3_218(.clk(clk),.reset(reset),.i1(intermediate_reg_2[77]),.i2(intermediate_reg_2[76]),.o(intermediate_reg_3[38])); 
mux_module mux_module_inst_3_219(.clk(clk),.reset(reset),.i1(intermediate_reg_2[75]),.i2(intermediate_reg_2[74]),.o(intermediate_reg_3[37]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_220(.clk(clk),.reset(reset),.i1(intermediate_reg_2[73]),.i2(intermediate_reg_2[72]),.o(intermediate_reg_3[36]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_221(.clk(clk),.reset(reset),.i1(intermediate_reg_2[71]),.i2(intermediate_reg_2[70]),.o(intermediate_reg_3[35])); 
fsm fsm_inst_3_222(.clk(clk),.reset(reset),.i1(intermediate_reg_2[69]),.i2(intermediate_reg_2[68]),.o(intermediate_reg_3[34])); 
mux_module mux_module_inst_3_223(.clk(clk),.reset(reset),.i1(intermediate_reg_2[67]),.i2(intermediate_reg_2[66]),.o(intermediate_reg_3[33]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_224(.clk(clk),.reset(reset),.i1(intermediate_reg_2[65]),.i2(intermediate_reg_2[64]),.o(intermediate_reg_3[32])); 
fsm fsm_inst_3_225(.clk(clk),.reset(reset),.i1(intermediate_reg_2[63]),.i2(intermediate_reg_2[62]),.o(intermediate_reg_3[31])); 
fsm fsm_inst_3_226(.clk(clk),.reset(reset),.i1(intermediate_reg_2[61]),.i2(intermediate_reg_2[60]),.o(intermediate_reg_3[30])); 
mux_module mux_module_inst_3_227(.clk(clk),.reset(reset),.i1(intermediate_reg_2[59]),.i2(intermediate_reg_2[58]),.o(intermediate_reg_3[29]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_228(.clk(clk),.reset(reset),.i1(intermediate_reg_2[57]),.i2(intermediate_reg_2[56]),.o(intermediate_reg_3[28]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_229(.clk(clk),.reset(reset),.i1(intermediate_reg_2[55]),.i2(intermediate_reg_2[54]),.o(intermediate_reg_3[27]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_230(.clk(clk),.reset(reset),.i1(intermediate_reg_2[53]),.i2(intermediate_reg_2[52]),.o(intermediate_reg_3[26])); 
mux_module mux_module_inst_3_231(.clk(clk),.reset(reset),.i1(intermediate_reg_2[51]),.i2(intermediate_reg_2[50]),.o(intermediate_reg_3[25]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_232(.clk(clk),.reset(reset),.i1(intermediate_reg_2[49]),.i2(intermediate_reg_2[48]),.o(intermediate_reg_3[24]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_233(.clk(clk),.reset(reset),.i1(intermediate_reg_2[47]),.i2(intermediate_reg_2[46]),.o(intermediate_reg_3[23])); 
mux_module mux_module_inst_3_234(.clk(clk),.reset(reset),.i1(intermediate_reg_2[45]),.i2(intermediate_reg_2[44]),.o(intermediate_reg_3[22]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_235(.clk(clk),.reset(reset),.i1(intermediate_reg_2[43]),.i2(intermediate_reg_2[42]),.o(intermediate_reg_3[21])); 
fsm fsm_inst_3_236(.clk(clk),.reset(reset),.i1(intermediate_reg_2[41]),.i2(intermediate_reg_2[40]),.o(intermediate_reg_3[20])); 
fsm fsm_inst_3_237(.clk(clk),.reset(reset),.i1(intermediate_reg_2[39]),.i2(intermediate_reg_2[38]),.o(intermediate_reg_3[19])); 
fsm fsm_inst_3_238(.clk(clk),.reset(reset),.i1(intermediate_reg_2[37]),.i2(intermediate_reg_2[36]),.o(intermediate_reg_3[18])); 
fsm fsm_inst_3_239(.clk(clk),.reset(reset),.i1(intermediate_reg_2[35]),.i2(intermediate_reg_2[34]),.o(intermediate_reg_3[17])); 
fsm fsm_inst_3_240(.clk(clk),.reset(reset),.i1(intermediate_reg_2[33]),.i2(intermediate_reg_2[32]),.o(intermediate_reg_3[16])); 
mux_module mux_module_inst_3_241(.clk(clk),.reset(reset),.i1(intermediate_reg_2[31]),.i2(intermediate_reg_2[30]),.o(intermediate_reg_3[15]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_242(.clk(clk),.reset(reset),.i1(intermediate_reg_2[29]),.i2(intermediate_reg_2[28]),.o(intermediate_reg_3[14]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_243(.clk(clk),.reset(reset),.i1(intermediate_reg_2[27]),.i2(intermediate_reg_2[26]),.o(intermediate_reg_3[13]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_244(.clk(clk),.reset(reset),.i1(intermediate_reg_2[25]),.i2(intermediate_reg_2[24]),.o(intermediate_reg_3[12])); 
fsm fsm_inst_3_245(.clk(clk),.reset(reset),.i1(intermediate_reg_2[23]),.i2(intermediate_reg_2[22]),.o(intermediate_reg_3[11])); 
fsm fsm_inst_3_246(.clk(clk),.reset(reset),.i1(intermediate_reg_2[21]),.i2(intermediate_reg_2[20]),.o(intermediate_reg_3[10])); 
fsm fsm_inst_3_247(.clk(clk),.reset(reset),.i1(intermediate_reg_2[19]),.i2(intermediate_reg_2[18]),.o(intermediate_reg_3[9])); 
fsm fsm_inst_3_248(.clk(clk),.reset(reset),.i1(intermediate_reg_2[17]),.i2(intermediate_reg_2[16]),.o(intermediate_reg_3[8])); 
fsm fsm_inst_3_249(.clk(clk),.reset(reset),.i1(intermediate_reg_2[15]),.i2(intermediate_reg_2[14]),.o(intermediate_reg_3[7])); 
fsm fsm_inst_3_250(.clk(clk),.reset(reset),.i1(intermediate_reg_2[13]),.i2(intermediate_reg_2[12]),.o(intermediate_reg_3[6])); 
fsm fsm_inst_3_251(.clk(clk),.reset(reset),.i1(intermediate_reg_2[11]),.i2(intermediate_reg_2[10]),.o(intermediate_reg_3[5])); 
fsm fsm_inst_3_252(.clk(clk),.reset(reset),.i1(intermediate_reg_2[9]),.i2(intermediate_reg_2[8]),.o(intermediate_reg_3[4])); 
mux_module mux_module_inst_3_253(.clk(clk),.reset(reset),.i1(intermediate_reg_2[7]),.i2(intermediate_reg_2[6]),.o(intermediate_reg_3[3]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_254(.clk(clk),.reset(reset),.i1(intermediate_reg_2[5]),.i2(intermediate_reg_2[4]),.o(intermediate_reg_3[2])); 
mux_module mux_module_inst_3_255(.clk(clk),.reset(reset),.i1(intermediate_reg_2[3]),.i2(intermediate_reg_2[2]),.o(intermediate_reg_3[1]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_256(.clk(clk),.reset(reset),.i1(intermediate_reg_2[1]),.i2(intermediate_reg_2[0]),.o(intermediate_reg_3[0])); 
wire [255:0]intermediate_wire_4; 
assign intermediate_wire_4[255] = intermediate_reg_3[256]^intermediate_reg_3[255] ; 
assign intermediate_wire_4[254:0] = intermediate_reg_3[254:0] ; 
always@(posedge clk) begin 
outp [255:0] <= intermediate_wire_4; 
outp[311:256] <= intermediate_wire_4[55:0] ; 
end 
endmodule 
 

module interface_23(input reg [9679:0] inp, output reg [9599:0] outp, input clk, input reset);
reg [9679:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [4839:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9679]),.i2(intermediate_reg_0[9678]),.o(intermediate_reg_1[4839]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9677]),.i2(intermediate_reg_0[9676]),.o(intermediate_reg_1[4838]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9675]),.i2(intermediate_reg_0[9674]),.o(intermediate_reg_1[4837]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9673]),.i2(intermediate_reg_0[9672]),.o(intermediate_reg_1[4836])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9671]),.i2(intermediate_reg_0[9670]),.o(intermediate_reg_1[4835]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9669]),.i2(intermediate_reg_0[9668]),.o(intermediate_reg_1[4834])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9667]),.i2(intermediate_reg_0[9666]),.o(intermediate_reg_1[4833]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9665]),.i2(intermediate_reg_0[9664]),.o(intermediate_reg_1[4832])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9663]),.i2(intermediate_reg_0[9662]),.o(intermediate_reg_1[4831]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9661]),.i2(intermediate_reg_0[9660]),.o(intermediate_reg_1[4830]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9659]),.i2(intermediate_reg_0[9658]),.o(intermediate_reg_1[4829])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9657]),.i2(intermediate_reg_0[9656]),.o(intermediate_reg_1[4828])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9655]),.i2(intermediate_reg_0[9654]),.o(intermediate_reg_1[4827]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9653]),.i2(intermediate_reg_0[9652]),.o(intermediate_reg_1[4826]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9651]),.i2(intermediate_reg_0[9650]),.o(intermediate_reg_1[4825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9649]),.i2(intermediate_reg_0[9648]),.o(intermediate_reg_1[4824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9647]),.i2(intermediate_reg_0[9646]),.o(intermediate_reg_1[4823]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9645]),.i2(intermediate_reg_0[9644]),.o(intermediate_reg_1[4822])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9643]),.i2(intermediate_reg_0[9642]),.o(intermediate_reg_1[4821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9641]),.i2(intermediate_reg_0[9640]),.o(intermediate_reg_1[4820]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9639]),.i2(intermediate_reg_0[9638]),.o(intermediate_reg_1[4819]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9637]),.i2(intermediate_reg_0[9636]),.o(intermediate_reg_1[4818])); 
fsm fsm_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9635]),.i2(intermediate_reg_0[9634]),.o(intermediate_reg_1[4817])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9633]),.i2(intermediate_reg_0[9632]),.o(intermediate_reg_1[4816]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9631]),.i2(intermediate_reg_0[9630]),.o(intermediate_reg_1[4815])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9629]),.i2(intermediate_reg_0[9628]),.o(intermediate_reg_1[4814]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9627]),.i2(intermediate_reg_0[9626]),.o(intermediate_reg_1[4813]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9625]),.i2(intermediate_reg_0[9624]),.o(intermediate_reg_1[4812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9623]),.i2(intermediate_reg_0[9622]),.o(intermediate_reg_1[4811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9621]),.i2(intermediate_reg_0[9620]),.o(intermediate_reg_1[4810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9619]),.i2(intermediate_reg_0[9618]),.o(intermediate_reg_1[4809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9617]),.i2(intermediate_reg_0[9616]),.o(intermediate_reg_1[4808]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9615]),.i2(intermediate_reg_0[9614]),.o(intermediate_reg_1[4807])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9613]),.i2(intermediate_reg_0[9612]),.o(intermediate_reg_1[4806]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9611]),.i2(intermediate_reg_0[9610]),.o(intermediate_reg_1[4805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9609]),.i2(intermediate_reg_0[9608]),.o(intermediate_reg_1[4804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9607]),.i2(intermediate_reg_0[9606]),.o(intermediate_reg_1[4803]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9605]),.i2(intermediate_reg_0[9604]),.o(intermediate_reg_1[4802])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9603]),.i2(intermediate_reg_0[9602]),.o(intermediate_reg_1[4801]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9601]),.i2(intermediate_reg_0[9600]),.o(intermediate_reg_1[4800]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9599]),.i2(intermediate_reg_0[9598]),.o(intermediate_reg_1[4799])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9597]),.i2(intermediate_reg_0[9596]),.o(intermediate_reg_1[4798])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9595]),.i2(intermediate_reg_0[9594]),.o(intermediate_reg_1[4797]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9593]),.i2(intermediate_reg_0[9592]),.o(intermediate_reg_1[4796])); 
fsm fsm_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9591]),.i2(intermediate_reg_0[9590]),.o(intermediate_reg_1[4795])); 
fsm fsm_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9589]),.i2(intermediate_reg_0[9588]),.o(intermediate_reg_1[4794])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9587]),.i2(intermediate_reg_0[9586]),.o(intermediate_reg_1[4793])); 
fsm fsm_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9585]),.i2(intermediate_reg_0[9584]),.o(intermediate_reg_1[4792])); 
fsm fsm_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9583]),.i2(intermediate_reg_0[9582]),.o(intermediate_reg_1[4791])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9581]),.i2(intermediate_reg_0[9580]),.o(intermediate_reg_1[4790]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9579]),.i2(intermediate_reg_0[9578]),.o(intermediate_reg_1[4789])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9577]),.i2(intermediate_reg_0[9576]),.o(intermediate_reg_1[4788]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9575]),.i2(intermediate_reg_0[9574]),.o(intermediate_reg_1[4787])); 
fsm fsm_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9573]),.i2(intermediate_reg_0[9572]),.o(intermediate_reg_1[4786])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9571]),.i2(intermediate_reg_0[9570]),.o(intermediate_reg_1[4785]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9569]),.i2(intermediate_reg_0[9568]),.o(intermediate_reg_1[4784])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9567]),.i2(intermediate_reg_0[9566]),.o(intermediate_reg_1[4783]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9565]),.i2(intermediate_reg_0[9564]),.o(intermediate_reg_1[4782])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9563]),.i2(intermediate_reg_0[9562]),.o(intermediate_reg_1[4781]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9561]),.i2(intermediate_reg_0[9560]),.o(intermediate_reg_1[4780]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9559]),.i2(intermediate_reg_0[9558]),.o(intermediate_reg_1[4779])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9557]),.i2(intermediate_reg_0[9556]),.o(intermediate_reg_1[4778]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9555]),.i2(intermediate_reg_0[9554]),.o(intermediate_reg_1[4777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9553]),.i2(intermediate_reg_0[9552]),.o(intermediate_reg_1[4776]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9551]),.i2(intermediate_reg_0[9550]),.o(intermediate_reg_1[4775])); 
fsm fsm_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9549]),.i2(intermediate_reg_0[9548]),.o(intermediate_reg_1[4774])); 
fsm fsm_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9547]),.i2(intermediate_reg_0[9546]),.o(intermediate_reg_1[4773])); 
fsm fsm_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9545]),.i2(intermediate_reg_0[9544]),.o(intermediate_reg_1[4772])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9543]),.i2(intermediate_reg_0[9542]),.o(intermediate_reg_1[4771]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9541]),.i2(intermediate_reg_0[9540]),.o(intermediate_reg_1[4770]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9539]),.i2(intermediate_reg_0[9538]),.o(intermediate_reg_1[4769])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9537]),.i2(intermediate_reg_0[9536]),.o(intermediate_reg_1[4768]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9535]),.i2(intermediate_reg_0[9534]),.o(intermediate_reg_1[4767])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9533]),.i2(intermediate_reg_0[9532]),.o(intermediate_reg_1[4766]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9531]),.i2(intermediate_reg_0[9530]),.o(intermediate_reg_1[4765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9529]),.i2(intermediate_reg_0[9528]),.o(intermediate_reg_1[4764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9527]),.i2(intermediate_reg_0[9526]),.o(intermediate_reg_1[4763]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9525]),.i2(intermediate_reg_0[9524]),.o(intermediate_reg_1[4762])); 
fsm fsm_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9523]),.i2(intermediate_reg_0[9522]),.o(intermediate_reg_1[4761])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9521]),.i2(intermediate_reg_0[9520]),.o(intermediate_reg_1[4760]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9519]),.i2(intermediate_reg_0[9518]),.o(intermediate_reg_1[4759])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9517]),.i2(intermediate_reg_0[9516]),.o(intermediate_reg_1[4758])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9515]),.i2(intermediate_reg_0[9514]),.o(intermediate_reg_1[4757]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9513]),.i2(intermediate_reg_0[9512]),.o(intermediate_reg_1[4756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9511]),.i2(intermediate_reg_0[9510]),.o(intermediate_reg_1[4755]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9509]),.i2(intermediate_reg_0[9508]),.o(intermediate_reg_1[4754])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9507]),.i2(intermediate_reg_0[9506]),.o(intermediate_reg_1[4753]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9505]),.i2(intermediate_reg_0[9504]),.o(intermediate_reg_1[4752])); 
fsm fsm_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9503]),.i2(intermediate_reg_0[9502]),.o(intermediate_reg_1[4751])); 
fsm fsm_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9501]),.i2(intermediate_reg_0[9500]),.o(intermediate_reg_1[4750])); 
fsm fsm_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9499]),.i2(intermediate_reg_0[9498]),.o(intermediate_reg_1[4749])); 
fsm fsm_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9497]),.i2(intermediate_reg_0[9496]),.o(intermediate_reg_1[4748])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9495]),.i2(intermediate_reg_0[9494]),.o(intermediate_reg_1[4747]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9493]),.i2(intermediate_reg_0[9492]),.o(intermediate_reg_1[4746])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9491]),.i2(intermediate_reg_0[9490]),.o(intermediate_reg_1[4745]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9489]),.i2(intermediate_reg_0[9488]),.o(intermediate_reg_1[4744])); 
fsm fsm_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9487]),.i2(intermediate_reg_0[9486]),.o(intermediate_reg_1[4743])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9485]),.i2(intermediate_reg_0[9484]),.o(intermediate_reg_1[4742]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9483]),.i2(intermediate_reg_0[9482]),.o(intermediate_reg_1[4741])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9481]),.i2(intermediate_reg_0[9480]),.o(intermediate_reg_1[4740]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9479]),.i2(intermediate_reg_0[9478]),.o(intermediate_reg_1[4739])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9477]),.i2(intermediate_reg_0[9476]),.o(intermediate_reg_1[4738])); 
fsm fsm_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9475]),.i2(intermediate_reg_0[9474]),.o(intermediate_reg_1[4737])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9473]),.i2(intermediate_reg_0[9472]),.o(intermediate_reg_1[4736]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9471]),.i2(intermediate_reg_0[9470]),.o(intermediate_reg_1[4735]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9469]),.i2(intermediate_reg_0[9468]),.o(intermediate_reg_1[4734])); 
fsm fsm_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9467]),.i2(intermediate_reg_0[9466]),.o(intermediate_reg_1[4733])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9465]),.i2(intermediate_reg_0[9464]),.o(intermediate_reg_1[4732]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9463]),.i2(intermediate_reg_0[9462]),.o(intermediate_reg_1[4731])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9461]),.i2(intermediate_reg_0[9460]),.o(intermediate_reg_1[4730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9459]),.i2(intermediate_reg_0[9458]),.o(intermediate_reg_1[4729]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9457]),.i2(intermediate_reg_0[9456]),.o(intermediate_reg_1[4728])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9455]),.i2(intermediate_reg_0[9454]),.o(intermediate_reg_1[4727])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9453]),.i2(intermediate_reg_0[9452]),.o(intermediate_reg_1[4726]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9451]),.i2(intermediate_reg_0[9450]),.o(intermediate_reg_1[4725])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9449]),.i2(intermediate_reg_0[9448]),.o(intermediate_reg_1[4724]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9447]),.i2(intermediate_reg_0[9446]),.o(intermediate_reg_1[4723])); 
fsm fsm_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9445]),.i2(intermediate_reg_0[9444]),.o(intermediate_reg_1[4722])); 
mux_module mux_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9443]),.i2(intermediate_reg_0[9442]),.o(intermediate_reg_1[4721]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9441]),.i2(intermediate_reg_0[9440]),.o(intermediate_reg_1[4720])); 
fsm fsm_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9439]),.i2(intermediate_reg_0[9438]),.o(intermediate_reg_1[4719])); 
fsm fsm_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9437]),.i2(intermediate_reg_0[9436]),.o(intermediate_reg_1[4718])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9435]),.i2(intermediate_reg_0[9434]),.o(intermediate_reg_1[4717]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9433]),.i2(intermediate_reg_0[9432]),.o(intermediate_reg_1[4716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9431]),.i2(intermediate_reg_0[9430]),.o(intermediate_reg_1[4715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9429]),.i2(intermediate_reg_0[9428]),.o(intermediate_reg_1[4714]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9427]),.i2(intermediate_reg_0[9426]),.o(intermediate_reg_1[4713]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9425]),.i2(intermediate_reg_0[9424]),.o(intermediate_reg_1[4712]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9423]),.i2(intermediate_reg_0[9422]),.o(intermediate_reg_1[4711])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9421]),.i2(intermediate_reg_0[9420]),.o(intermediate_reg_1[4710]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9419]),.i2(intermediate_reg_0[9418]),.o(intermediate_reg_1[4709])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9417]),.i2(intermediate_reg_0[9416]),.o(intermediate_reg_1[4708])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9415]),.i2(intermediate_reg_0[9414]),.o(intermediate_reg_1[4707]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9413]),.i2(intermediate_reg_0[9412]),.o(intermediate_reg_1[4706])); 
fsm fsm_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9411]),.i2(intermediate_reg_0[9410]),.o(intermediate_reg_1[4705])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9409]),.i2(intermediate_reg_0[9408]),.o(intermediate_reg_1[4704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9407]),.i2(intermediate_reg_0[9406]),.o(intermediate_reg_1[4703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9405]),.i2(intermediate_reg_0[9404]),.o(intermediate_reg_1[4702]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9403]),.i2(intermediate_reg_0[9402]),.o(intermediate_reg_1[4701])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9401]),.i2(intermediate_reg_0[9400]),.o(intermediate_reg_1[4700])); 
fsm fsm_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9399]),.i2(intermediate_reg_0[9398]),.o(intermediate_reg_1[4699])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9397]),.i2(intermediate_reg_0[9396]),.o(intermediate_reg_1[4698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9395]),.i2(intermediate_reg_0[9394]),.o(intermediate_reg_1[4697]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9393]),.i2(intermediate_reg_0[9392]),.o(intermediate_reg_1[4696])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9391]),.i2(intermediate_reg_0[9390]),.o(intermediate_reg_1[4695]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9389]),.i2(intermediate_reg_0[9388]),.o(intermediate_reg_1[4694])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9387]),.i2(intermediate_reg_0[9386]),.o(intermediate_reg_1[4693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9385]),.i2(intermediate_reg_0[9384]),.o(intermediate_reg_1[4692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9383]),.i2(intermediate_reg_0[9382]),.o(intermediate_reg_1[4691]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9381]),.i2(intermediate_reg_0[9380]),.o(intermediate_reg_1[4690]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9379]),.i2(intermediate_reg_0[9378]),.o(intermediate_reg_1[4689]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9377]),.i2(intermediate_reg_0[9376]),.o(intermediate_reg_1[4688])); 
fsm fsm_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9375]),.i2(intermediate_reg_0[9374]),.o(intermediate_reg_1[4687])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9373]),.i2(intermediate_reg_0[9372]),.o(intermediate_reg_1[4686])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9371]),.i2(intermediate_reg_0[9370]),.o(intermediate_reg_1[4685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9369]),.i2(intermediate_reg_0[9368]),.o(intermediate_reg_1[4684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9367]),.i2(intermediate_reg_0[9366]),.o(intermediate_reg_1[4683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9365]),.i2(intermediate_reg_0[9364]),.o(intermediate_reg_1[4682]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9363]),.i2(intermediate_reg_0[9362]),.o(intermediate_reg_1[4681])); 
mux_module mux_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9361]),.i2(intermediate_reg_0[9360]),.o(intermediate_reg_1[4680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9359]),.i2(intermediate_reg_0[9358]),.o(intermediate_reg_1[4679]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9357]),.i2(intermediate_reg_0[9356]),.o(intermediate_reg_1[4678])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9355]),.i2(intermediate_reg_0[9354]),.o(intermediate_reg_1[4677]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9353]),.i2(intermediate_reg_0[9352]),.o(intermediate_reg_1[4676])); 
mux_module mux_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9351]),.i2(intermediate_reg_0[9350]),.o(intermediate_reg_1[4675]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9349]),.i2(intermediate_reg_0[9348]),.o(intermediate_reg_1[4674])); 
mux_module mux_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9347]),.i2(intermediate_reg_0[9346]),.o(intermediate_reg_1[4673]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9345]),.i2(intermediate_reg_0[9344]),.o(intermediate_reg_1[4672])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9343]),.i2(intermediate_reg_0[9342]),.o(intermediate_reg_1[4671]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9341]),.i2(intermediate_reg_0[9340]),.o(intermediate_reg_1[4670])); 
fsm fsm_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9339]),.i2(intermediate_reg_0[9338]),.o(intermediate_reg_1[4669])); 
fsm fsm_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9337]),.i2(intermediate_reg_0[9336]),.o(intermediate_reg_1[4668])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9335]),.i2(intermediate_reg_0[9334]),.o(intermediate_reg_1[4667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9333]),.i2(intermediate_reg_0[9332]),.o(intermediate_reg_1[4666]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9331]),.i2(intermediate_reg_0[9330]),.o(intermediate_reg_1[4665])); 
fsm fsm_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9329]),.i2(intermediate_reg_0[9328]),.o(intermediate_reg_1[4664])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9327]),.i2(intermediate_reg_0[9326]),.o(intermediate_reg_1[4663])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9325]),.i2(intermediate_reg_0[9324]),.o(intermediate_reg_1[4662]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9323]),.i2(intermediate_reg_0[9322]),.o(intermediate_reg_1[4661])); 
fsm fsm_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9321]),.i2(intermediate_reg_0[9320]),.o(intermediate_reg_1[4660])); 
fsm fsm_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9319]),.i2(intermediate_reg_0[9318]),.o(intermediate_reg_1[4659])); 
fsm fsm_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9317]),.i2(intermediate_reg_0[9316]),.o(intermediate_reg_1[4658])); 
fsm fsm_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9315]),.i2(intermediate_reg_0[9314]),.o(intermediate_reg_1[4657])); 
fsm fsm_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9313]),.i2(intermediate_reg_0[9312]),.o(intermediate_reg_1[4656])); 
fsm fsm_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9311]),.i2(intermediate_reg_0[9310]),.o(intermediate_reg_1[4655])); 
fsm fsm_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9309]),.i2(intermediate_reg_0[9308]),.o(intermediate_reg_1[4654])); 
fsm fsm_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9307]),.i2(intermediate_reg_0[9306]),.o(intermediate_reg_1[4653])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9305]),.i2(intermediate_reg_0[9304]),.o(intermediate_reg_1[4652]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9303]),.i2(intermediate_reg_0[9302]),.o(intermediate_reg_1[4651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9301]),.i2(intermediate_reg_0[9300]),.o(intermediate_reg_1[4650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9299]),.i2(intermediate_reg_0[9298]),.o(intermediate_reg_1[4649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9297]),.i2(intermediate_reg_0[9296]),.o(intermediate_reg_1[4648]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9295]),.i2(intermediate_reg_0[9294]),.o(intermediate_reg_1[4647])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9293]),.i2(intermediate_reg_0[9292]),.o(intermediate_reg_1[4646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9291]),.i2(intermediate_reg_0[9290]),.o(intermediate_reg_1[4645]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9289]),.i2(intermediate_reg_0[9288]),.o(intermediate_reg_1[4644]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9287]),.i2(intermediate_reg_0[9286]),.o(intermediate_reg_1[4643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9285]),.i2(intermediate_reg_0[9284]),.o(intermediate_reg_1[4642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9283]),.i2(intermediate_reg_0[9282]),.o(intermediate_reg_1[4641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9281]),.i2(intermediate_reg_0[9280]),.o(intermediate_reg_1[4640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9279]),.i2(intermediate_reg_0[9278]),.o(intermediate_reg_1[4639]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9277]),.i2(intermediate_reg_0[9276]),.o(intermediate_reg_1[4638])); 
mux_module mux_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9275]),.i2(intermediate_reg_0[9274]),.o(intermediate_reg_1[4637]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9273]),.i2(intermediate_reg_0[9272]),.o(intermediate_reg_1[4636])); 
fsm fsm_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9271]),.i2(intermediate_reg_0[9270]),.o(intermediate_reg_1[4635])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9269]),.i2(intermediate_reg_0[9268]),.o(intermediate_reg_1[4634]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9267]),.i2(intermediate_reg_0[9266]),.o(intermediate_reg_1[4633])); 
mux_module mux_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9265]),.i2(intermediate_reg_0[9264]),.o(intermediate_reg_1[4632]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9263]),.i2(intermediate_reg_0[9262]),.o(intermediate_reg_1[4631]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9261]),.i2(intermediate_reg_0[9260]),.o(intermediate_reg_1[4630])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9259]),.i2(intermediate_reg_0[9258]),.o(intermediate_reg_1[4629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9257]),.i2(intermediate_reg_0[9256]),.o(intermediate_reg_1[4628]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9255]),.i2(intermediate_reg_0[9254]),.o(intermediate_reg_1[4627]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9253]),.i2(intermediate_reg_0[9252]),.o(intermediate_reg_1[4626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9251]),.i2(intermediate_reg_0[9250]),.o(intermediate_reg_1[4625])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9249]),.i2(intermediate_reg_0[9248]),.o(intermediate_reg_1[4624])); 
fsm fsm_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9247]),.i2(intermediate_reg_0[9246]),.o(intermediate_reg_1[4623])); 
mux_module mux_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9245]),.i2(intermediate_reg_0[9244]),.o(intermediate_reg_1[4622]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9243]),.i2(intermediate_reg_0[9242]),.o(intermediate_reg_1[4621]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9241]),.i2(intermediate_reg_0[9240]),.o(intermediate_reg_1[4620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9239]),.i2(intermediate_reg_0[9238]),.o(intermediate_reg_1[4619]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9237]),.i2(intermediate_reg_0[9236]),.o(intermediate_reg_1[4618])); 
fsm fsm_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9235]),.i2(intermediate_reg_0[9234]),.o(intermediate_reg_1[4617])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9233]),.i2(intermediate_reg_0[9232]),.o(intermediate_reg_1[4616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9231]),.i2(intermediate_reg_0[9230]),.o(intermediate_reg_1[4615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9229]),.i2(intermediate_reg_0[9228]),.o(intermediate_reg_1[4614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9227]),.i2(intermediate_reg_0[9226]),.o(intermediate_reg_1[4613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9225]),.i2(intermediate_reg_0[9224]),.o(intermediate_reg_1[4612]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9223]),.i2(intermediate_reg_0[9222]),.o(intermediate_reg_1[4611]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9221]),.i2(intermediate_reg_0[9220]),.o(intermediate_reg_1[4610]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9219]),.i2(intermediate_reg_0[9218]),.o(intermediate_reg_1[4609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9217]),.i2(intermediate_reg_0[9216]),.o(intermediate_reg_1[4608]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9215]),.i2(intermediate_reg_0[9214]),.o(intermediate_reg_1[4607])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9213]),.i2(intermediate_reg_0[9212]),.o(intermediate_reg_1[4606]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9211]),.i2(intermediate_reg_0[9210]),.o(intermediate_reg_1[4605])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9209]),.i2(intermediate_reg_0[9208]),.o(intermediate_reg_1[4604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9207]),.i2(intermediate_reg_0[9206]),.o(intermediate_reg_1[4603]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9205]),.i2(intermediate_reg_0[9204]),.o(intermediate_reg_1[4602])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9203]),.i2(intermediate_reg_0[9202]),.o(intermediate_reg_1[4601]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9201]),.i2(intermediate_reg_0[9200]),.o(intermediate_reg_1[4600]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9199]),.i2(intermediate_reg_0[9198]),.o(intermediate_reg_1[4599])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9197]),.i2(intermediate_reg_0[9196]),.o(intermediate_reg_1[4598])); 
fsm fsm_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9195]),.i2(intermediate_reg_0[9194]),.o(intermediate_reg_1[4597])); 
fsm fsm_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9193]),.i2(intermediate_reg_0[9192]),.o(intermediate_reg_1[4596])); 
fsm fsm_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9191]),.i2(intermediate_reg_0[9190]),.o(intermediate_reg_1[4595])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9189]),.i2(intermediate_reg_0[9188]),.o(intermediate_reg_1[4594])); 
fsm fsm_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9187]),.i2(intermediate_reg_0[9186]),.o(intermediate_reg_1[4593])); 
mux_module mux_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9185]),.i2(intermediate_reg_0[9184]),.o(intermediate_reg_1[4592]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9183]),.i2(intermediate_reg_0[9182]),.o(intermediate_reg_1[4591])); 
fsm fsm_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9181]),.i2(intermediate_reg_0[9180]),.o(intermediate_reg_1[4590])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9179]),.i2(intermediate_reg_0[9178]),.o(intermediate_reg_1[4589]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9177]),.i2(intermediate_reg_0[9176]),.o(intermediate_reg_1[4588])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9175]),.i2(intermediate_reg_0[9174]),.o(intermediate_reg_1[4587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9173]),.i2(intermediate_reg_0[9172]),.o(intermediate_reg_1[4586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9171]),.i2(intermediate_reg_0[9170]),.o(intermediate_reg_1[4585]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9169]),.i2(intermediate_reg_0[9168]),.o(intermediate_reg_1[4584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9167]),.i2(intermediate_reg_0[9166]),.o(intermediate_reg_1[4583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9165]),.i2(intermediate_reg_0[9164]),.o(intermediate_reg_1[4582]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9163]),.i2(intermediate_reg_0[9162]),.o(intermediate_reg_1[4581])); 
fsm fsm_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9161]),.i2(intermediate_reg_0[9160]),.o(intermediate_reg_1[4580])); 
fsm fsm_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9159]),.i2(intermediate_reg_0[9158]),.o(intermediate_reg_1[4579])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9157]),.i2(intermediate_reg_0[9156]),.o(intermediate_reg_1[4578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9155]),.i2(intermediate_reg_0[9154]),.o(intermediate_reg_1[4577]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9153]),.i2(intermediate_reg_0[9152]),.o(intermediate_reg_1[4576])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9151]),.i2(intermediate_reg_0[9150]),.o(intermediate_reg_1[4575]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9149]),.i2(intermediate_reg_0[9148]),.o(intermediate_reg_1[4574])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9147]),.i2(intermediate_reg_0[9146]),.o(intermediate_reg_1[4573]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9145]),.i2(intermediate_reg_0[9144]),.o(intermediate_reg_1[4572]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9143]),.i2(intermediate_reg_0[9142]),.o(intermediate_reg_1[4571])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9141]),.i2(intermediate_reg_0[9140]),.o(intermediate_reg_1[4570])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9139]),.i2(intermediate_reg_0[9138]),.o(intermediate_reg_1[4569]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9137]),.i2(intermediate_reg_0[9136]),.o(intermediate_reg_1[4568])); 
fsm fsm_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9135]),.i2(intermediate_reg_0[9134]),.o(intermediate_reg_1[4567])); 
mux_module mux_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9133]),.i2(intermediate_reg_0[9132]),.o(intermediate_reg_1[4566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9131]),.i2(intermediate_reg_0[9130]),.o(intermediate_reg_1[4565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9129]),.i2(intermediate_reg_0[9128]),.o(intermediate_reg_1[4564]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9127]),.i2(intermediate_reg_0[9126]),.o(intermediate_reg_1[4563])); 
fsm fsm_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9125]),.i2(intermediate_reg_0[9124]),.o(intermediate_reg_1[4562])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9123]),.i2(intermediate_reg_0[9122]),.o(intermediate_reg_1[4561]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9121]),.i2(intermediate_reg_0[9120]),.o(intermediate_reg_1[4560])); 
fsm fsm_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9119]),.i2(intermediate_reg_0[9118]),.o(intermediate_reg_1[4559])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9117]),.i2(intermediate_reg_0[9116]),.o(intermediate_reg_1[4558]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9115]),.i2(intermediate_reg_0[9114]),.o(intermediate_reg_1[4557])); 
mux_module mux_module_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9113]),.i2(intermediate_reg_0[9112]),.o(intermediate_reg_1[4556]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9111]),.i2(intermediate_reg_0[9110]),.o(intermediate_reg_1[4555]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9109]),.i2(intermediate_reg_0[9108]),.o(intermediate_reg_1[4554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9107]),.i2(intermediate_reg_0[9106]),.o(intermediate_reg_1[4553]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9105]),.i2(intermediate_reg_0[9104]),.o(intermediate_reg_1[4552])); 
fsm fsm_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9103]),.i2(intermediate_reg_0[9102]),.o(intermediate_reg_1[4551])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9101]),.i2(intermediate_reg_0[9100]),.o(intermediate_reg_1[4550]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9099]),.i2(intermediate_reg_0[9098]),.o(intermediate_reg_1[4549])); 
mux_module mux_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9097]),.i2(intermediate_reg_0[9096]),.o(intermediate_reg_1[4548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9095]),.i2(intermediate_reg_0[9094]),.o(intermediate_reg_1[4547]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9093]),.i2(intermediate_reg_0[9092]),.o(intermediate_reg_1[4546])); 
fsm fsm_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9091]),.i2(intermediate_reg_0[9090]),.o(intermediate_reg_1[4545])); 
mux_module mux_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9089]),.i2(intermediate_reg_0[9088]),.o(intermediate_reg_1[4544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9087]),.i2(intermediate_reg_0[9086]),.o(intermediate_reg_1[4543]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9085]),.i2(intermediate_reg_0[9084]),.o(intermediate_reg_1[4542])); 
fsm fsm_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9083]),.i2(intermediate_reg_0[9082]),.o(intermediate_reg_1[4541])); 
mux_module mux_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9081]),.i2(intermediate_reg_0[9080]),.o(intermediate_reg_1[4540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9079]),.i2(intermediate_reg_0[9078]),.o(intermediate_reg_1[4539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9077]),.i2(intermediate_reg_0[9076]),.o(intermediate_reg_1[4538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9075]),.i2(intermediate_reg_0[9074]),.o(intermediate_reg_1[4537]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9073]),.i2(intermediate_reg_0[9072]),.o(intermediate_reg_1[4536])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9071]),.i2(intermediate_reg_0[9070]),.o(intermediate_reg_1[4535])); 
fsm fsm_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9069]),.i2(intermediate_reg_0[9068]),.o(intermediate_reg_1[4534])); 
fsm fsm_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9067]),.i2(intermediate_reg_0[9066]),.o(intermediate_reg_1[4533])); 
fsm fsm_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9065]),.i2(intermediate_reg_0[9064]),.o(intermediate_reg_1[4532])); 
fsm fsm_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9063]),.i2(intermediate_reg_0[9062]),.o(intermediate_reg_1[4531])); 
fsm fsm_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9061]),.i2(intermediate_reg_0[9060]),.o(intermediate_reg_1[4530])); 
mux_module mux_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9059]),.i2(intermediate_reg_0[9058]),.o(intermediate_reg_1[4529]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9057]),.i2(intermediate_reg_0[9056]),.o(intermediate_reg_1[4528])); 
fsm fsm_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9055]),.i2(intermediate_reg_0[9054]),.o(intermediate_reg_1[4527])); 
mux_module mux_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9053]),.i2(intermediate_reg_0[9052]),.o(intermediate_reg_1[4526]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9051]),.i2(intermediate_reg_0[9050]),.o(intermediate_reg_1[4525])); 
fsm fsm_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9049]),.i2(intermediate_reg_0[9048]),.o(intermediate_reg_1[4524])); 
fsm fsm_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9047]),.i2(intermediate_reg_0[9046]),.o(intermediate_reg_1[4523])); 
fsm fsm_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9045]),.i2(intermediate_reg_0[9044]),.o(intermediate_reg_1[4522])); 
fsm fsm_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9043]),.i2(intermediate_reg_0[9042]),.o(intermediate_reg_1[4521])); 
fsm fsm_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9041]),.i2(intermediate_reg_0[9040]),.o(intermediate_reg_1[4520])); 
fsm fsm_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9039]),.i2(intermediate_reg_0[9038]),.o(intermediate_reg_1[4519])); 
fsm fsm_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9037]),.i2(intermediate_reg_0[9036]),.o(intermediate_reg_1[4518])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9035]),.i2(intermediate_reg_0[9034]),.o(intermediate_reg_1[4517])); 
fsm fsm_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9033]),.i2(intermediate_reg_0[9032]),.o(intermediate_reg_1[4516])); 
mux_module mux_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9031]),.i2(intermediate_reg_0[9030]),.o(intermediate_reg_1[4515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9029]),.i2(intermediate_reg_0[9028]),.o(intermediate_reg_1[4514]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9027]),.i2(intermediate_reg_0[9026]),.o(intermediate_reg_1[4513])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9025]),.i2(intermediate_reg_0[9024]),.o(intermediate_reg_1[4512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9023]),.i2(intermediate_reg_0[9022]),.o(intermediate_reg_1[4511]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9021]),.i2(intermediate_reg_0[9020]),.o(intermediate_reg_1[4510])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9019]),.i2(intermediate_reg_0[9018]),.o(intermediate_reg_1[4509]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9017]),.i2(intermediate_reg_0[9016]),.o(intermediate_reg_1[4508])); 
mux_module mux_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9015]),.i2(intermediate_reg_0[9014]),.o(intermediate_reg_1[4507]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9013]),.i2(intermediate_reg_0[9012]),.o(intermediate_reg_1[4506])); 
fsm fsm_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9011]),.i2(intermediate_reg_0[9010]),.o(intermediate_reg_1[4505])); 
fsm fsm_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9009]),.i2(intermediate_reg_0[9008]),.o(intermediate_reg_1[4504])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9007]),.i2(intermediate_reg_0[9006]),.o(intermediate_reg_1[4503]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9005]),.i2(intermediate_reg_0[9004]),.o(intermediate_reg_1[4502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9003]),.i2(intermediate_reg_0[9002]),.o(intermediate_reg_1[4501]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9001]),.i2(intermediate_reg_0[9000]),.o(intermediate_reg_1[4500])); 
fsm fsm_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8999]),.i2(intermediate_reg_0[8998]),.o(intermediate_reg_1[4499])); 
fsm fsm_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8997]),.i2(intermediate_reg_0[8996]),.o(intermediate_reg_1[4498])); 
fsm fsm_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8995]),.i2(intermediate_reg_0[8994]),.o(intermediate_reg_1[4497])); 
fsm fsm_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8993]),.i2(intermediate_reg_0[8992]),.o(intermediate_reg_1[4496])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8991]),.i2(intermediate_reg_0[8990]),.o(intermediate_reg_1[4495])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8989]),.i2(intermediate_reg_0[8988]),.o(intermediate_reg_1[4494])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8987]),.i2(intermediate_reg_0[8986]),.o(intermediate_reg_1[4493])); 
fsm fsm_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8985]),.i2(intermediate_reg_0[8984]),.o(intermediate_reg_1[4492])); 
fsm fsm_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8983]),.i2(intermediate_reg_0[8982]),.o(intermediate_reg_1[4491])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8981]),.i2(intermediate_reg_0[8980]),.o(intermediate_reg_1[4490]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8979]),.i2(intermediate_reg_0[8978]),.o(intermediate_reg_1[4489])); 
mux_module mux_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8977]),.i2(intermediate_reg_0[8976]),.o(intermediate_reg_1[4488]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8975]),.i2(intermediate_reg_0[8974]),.o(intermediate_reg_1[4487])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8973]),.i2(intermediate_reg_0[8972]),.o(intermediate_reg_1[4486]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8971]),.i2(intermediate_reg_0[8970]),.o(intermediate_reg_1[4485])); 
mux_module mux_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8969]),.i2(intermediate_reg_0[8968]),.o(intermediate_reg_1[4484]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8967]),.i2(intermediate_reg_0[8966]),.o(intermediate_reg_1[4483])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8965]),.i2(intermediate_reg_0[8964]),.o(intermediate_reg_1[4482]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8963]),.i2(intermediate_reg_0[8962]),.o(intermediate_reg_1[4481])); 
fsm fsm_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8961]),.i2(intermediate_reg_0[8960]),.o(intermediate_reg_1[4480])); 
fsm fsm_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8959]),.i2(intermediate_reg_0[8958]),.o(intermediate_reg_1[4479])); 
mux_module mux_module_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8957]),.i2(intermediate_reg_0[8956]),.o(intermediate_reg_1[4478]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8955]),.i2(intermediate_reg_0[8954]),.o(intermediate_reg_1[4477]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8953]),.i2(intermediate_reg_0[8952]),.o(intermediate_reg_1[4476])); 
mux_module mux_module_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8951]),.i2(intermediate_reg_0[8950]),.o(intermediate_reg_1[4475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8949]),.i2(intermediate_reg_0[8948]),.o(intermediate_reg_1[4474]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8947]),.i2(intermediate_reg_0[8946]),.o(intermediate_reg_1[4473])); 
fsm fsm_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8945]),.i2(intermediate_reg_0[8944]),.o(intermediate_reg_1[4472])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8943]),.i2(intermediate_reg_0[8942]),.o(intermediate_reg_1[4471]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8941]),.i2(intermediate_reg_0[8940]),.o(intermediate_reg_1[4470]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8939]),.i2(intermediate_reg_0[8938]),.o(intermediate_reg_1[4469])); 
fsm fsm_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8937]),.i2(intermediate_reg_0[8936]),.o(intermediate_reg_1[4468])); 
fsm fsm_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8935]),.i2(intermediate_reg_0[8934]),.o(intermediate_reg_1[4467])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8933]),.i2(intermediate_reg_0[8932]),.o(intermediate_reg_1[4466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8931]),.i2(intermediate_reg_0[8930]),.o(intermediate_reg_1[4465]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8929]),.i2(intermediate_reg_0[8928]),.o(intermediate_reg_1[4464])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8927]),.i2(intermediate_reg_0[8926]),.o(intermediate_reg_1[4463])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8925]),.i2(intermediate_reg_0[8924]),.o(intermediate_reg_1[4462]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8923]),.i2(intermediate_reg_0[8922]),.o(intermediate_reg_1[4461])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8921]),.i2(intermediate_reg_0[8920]),.o(intermediate_reg_1[4460])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8919]),.i2(intermediate_reg_0[8918]),.o(intermediate_reg_1[4459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8917]),.i2(intermediate_reg_0[8916]),.o(intermediate_reg_1[4458]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8915]),.i2(intermediate_reg_0[8914]),.o(intermediate_reg_1[4457])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8913]),.i2(intermediate_reg_0[8912]),.o(intermediate_reg_1[4456]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8911]),.i2(intermediate_reg_0[8910]),.o(intermediate_reg_1[4455])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8909]),.i2(intermediate_reg_0[8908]),.o(intermediate_reg_1[4454]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8907]),.i2(intermediate_reg_0[8906]),.o(intermediate_reg_1[4453])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8905]),.i2(intermediate_reg_0[8904]),.o(intermediate_reg_1[4452]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8903]),.i2(intermediate_reg_0[8902]),.o(intermediate_reg_1[4451])); 
fsm fsm_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8901]),.i2(intermediate_reg_0[8900]),.o(intermediate_reg_1[4450])); 
fsm fsm_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8899]),.i2(intermediate_reg_0[8898]),.o(intermediate_reg_1[4449])); 
fsm fsm_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8897]),.i2(intermediate_reg_0[8896]),.o(intermediate_reg_1[4448])); 
mux_module mux_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8895]),.i2(intermediate_reg_0[8894]),.o(intermediate_reg_1[4447]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8893]),.i2(intermediate_reg_0[8892]),.o(intermediate_reg_1[4446])); 
fsm fsm_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8891]),.i2(intermediate_reg_0[8890]),.o(intermediate_reg_1[4445])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8889]),.i2(intermediate_reg_0[8888]),.o(intermediate_reg_1[4444])); 
fsm fsm_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8887]),.i2(intermediate_reg_0[8886]),.o(intermediate_reg_1[4443])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8885]),.i2(intermediate_reg_0[8884]),.o(intermediate_reg_1[4442])); 
mux_module mux_module_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8883]),.i2(intermediate_reg_0[8882]),.o(intermediate_reg_1[4441]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8881]),.i2(intermediate_reg_0[8880]),.o(intermediate_reg_1[4440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8879]),.i2(intermediate_reg_0[8878]),.o(intermediate_reg_1[4439]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8877]),.i2(intermediate_reg_0[8876]),.o(intermediate_reg_1[4438])); 
mux_module mux_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8875]),.i2(intermediate_reg_0[8874]),.o(intermediate_reg_1[4437]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8873]),.i2(intermediate_reg_0[8872]),.o(intermediate_reg_1[4436])); 
fsm fsm_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8871]),.i2(intermediate_reg_0[8870]),.o(intermediate_reg_1[4435])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8869]),.i2(intermediate_reg_0[8868]),.o(intermediate_reg_1[4434])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8867]),.i2(intermediate_reg_0[8866]),.o(intermediate_reg_1[4433])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8865]),.i2(intermediate_reg_0[8864]),.o(intermediate_reg_1[4432])); 
fsm fsm_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8863]),.i2(intermediate_reg_0[8862]),.o(intermediate_reg_1[4431])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8861]),.i2(intermediate_reg_0[8860]),.o(intermediate_reg_1[4430]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8859]),.i2(intermediate_reg_0[8858]),.o(intermediate_reg_1[4429])); 
fsm fsm_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8857]),.i2(intermediate_reg_0[8856]),.o(intermediate_reg_1[4428])); 
fsm fsm_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8855]),.i2(intermediate_reg_0[8854]),.o(intermediate_reg_1[4427])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8853]),.i2(intermediate_reg_0[8852]),.o(intermediate_reg_1[4426])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8851]),.i2(intermediate_reg_0[8850]),.o(intermediate_reg_1[4425]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8849]),.i2(intermediate_reg_0[8848]),.o(intermediate_reg_1[4424])); 
fsm fsm_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8847]),.i2(intermediate_reg_0[8846]),.o(intermediate_reg_1[4423])); 
mux_module mux_module_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8845]),.i2(intermediate_reg_0[8844]),.o(intermediate_reg_1[4422]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8843]),.i2(intermediate_reg_0[8842]),.o(intermediate_reg_1[4421]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8841]),.i2(intermediate_reg_0[8840]),.o(intermediate_reg_1[4420]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8839]),.i2(intermediate_reg_0[8838]),.o(intermediate_reg_1[4419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8837]),.i2(intermediate_reg_0[8836]),.o(intermediate_reg_1[4418]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8835]),.i2(intermediate_reg_0[8834]),.o(intermediate_reg_1[4417])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8833]),.i2(intermediate_reg_0[8832]),.o(intermediate_reg_1[4416])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8831]),.i2(intermediate_reg_0[8830]),.o(intermediate_reg_1[4415])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8829]),.i2(intermediate_reg_0[8828]),.o(intermediate_reg_1[4414])); 
mux_module mux_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8827]),.i2(intermediate_reg_0[8826]),.o(intermediate_reg_1[4413]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8825]),.i2(intermediate_reg_0[8824]),.o(intermediate_reg_1[4412])); 
fsm fsm_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8823]),.i2(intermediate_reg_0[8822]),.o(intermediate_reg_1[4411])); 
fsm fsm_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8821]),.i2(intermediate_reg_0[8820]),.o(intermediate_reg_1[4410])); 
fsm fsm_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8819]),.i2(intermediate_reg_0[8818]),.o(intermediate_reg_1[4409])); 
fsm fsm_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8817]),.i2(intermediate_reg_0[8816]),.o(intermediate_reg_1[4408])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8815]),.i2(intermediate_reg_0[8814]),.o(intermediate_reg_1[4407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8813]),.i2(intermediate_reg_0[8812]),.o(intermediate_reg_1[4406])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8811]),.i2(intermediate_reg_0[8810]),.o(intermediate_reg_1[4405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8809]),.i2(intermediate_reg_0[8808]),.o(intermediate_reg_1[4404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8807]),.i2(intermediate_reg_0[8806]),.o(intermediate_reg_1[4403])); 
mux_module mux_module_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8805]),.i2(intermediate_reg_0[8804]),.o(intermediate_reg_1[4402]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8803]),.i2(intermediate_reg_0[8802]),.o(intermediate_reg_1[4401]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8801]),.i2(intermediate_reg_0[8800]),.o(intermediate_reg_1[4400]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8799]),.i2(intermediate_reg_0[8798]),.o(intermediate_reg_1[4399])); 
mux_module mux_module_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8797]),.i2(intermediate_reg_0[8796]),.o(intermediate_reg_1[4398]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8795]),.i2(intermediate_reg_0[8794]),.o(intermediate_reg_1[4397])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8793]),.i2(intermediate_reg_0[8792]),.o(intermediate_reg_1[4396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8791]),.i2(intermediate_reg_0[8790]),.o(intermediate_reg_1[4395]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8789]),.i2(intermediate_reg_0[8788]),.o(intermediate_reg_1[4394])); 
mux_module mux_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8787]),.i2(intermediate_reg_0[8786]),.o(intermediate_reg_1[4393]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8785]),.i2(intermediate_reg_0[8784]),.o(intermediate_reg_1[4392]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8783]),.i2(intermediate_reg_0[8782]),.o(intermediate_reg_1[4391]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8781]),.i2(intermediate_reg_0[8780]),.o(intermediate_reg_1[4390]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8779]),.i2(intermediate_reg_0[8778]),.o(intermediate_reg_1[4389]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8777]),.i2(intermediate_reg_0[8776]),.o(intermediate_reg_1[4388])); 
fsm fsm_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8775]),.i2(intermediate_reg_0[8774]),.o(intermediate_reg_1[4387])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8773]),.i2(intermediate_reg_0[8772]),.o(intermediate_reg_1[4386])); 
mux_module mux_module_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8771]),.i2(intermediate_reg_0[8770]),.o(intermediate_reg_1[4385]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8769]),.i2(intermediate_reg_0[8768]),.o(intermediate_reg_1[4384])); 
fsm fsm_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8767]),.i2(intermediate_reg_0[8766]),.o(intermediate_reg_1[4383])); 
fsm fsm_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8765]),.i2(intermediate_reg_0[8764]),.o(intermediate_reg_1[4382])); 
mux_module mux_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8763]),.i2(intermediate_reg_0[8762]),.o(intermediate_reg_1[4381]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8761]),.i2(intermediate_reg_0[8760]),.o(intermediate_reg_1[4380]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8759]),.i2(intermediate_reg_0[8758]),.o(intermediate_reg_1[4379])); 
mux_module mux_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8757]),.i2(intermediate_reg_0[8756]),.o(intermediate_reg_1[4378]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8755]),.i2(intermediate_reg_0[8754]),.o(intermediate_reg_1[4377])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8753]),.i2(intermediate_reg_0[8752]),.o(intermediate_reg_1[4376]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8751]),.i2(intermediate_reg_0[8750]),.o(intermediate_reg_1[4375]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8749]),.i2(intermediate_reg_0[8748]),.o(intermediate_reg_1[4374])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8747]),.i2(intermediate_reg_0[8746]),.o(intermediate_reg_1[4373])); 
mux_module mux_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8745]),.i2(intermediate_reg_0[8744]),.o(intermediate_reg_1[4372]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8743]),.i2(intermediate_reg_0[8742]),.o(intermediate_reg_1[4371])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8741]),.i2(intermediate_reg_0[8740]),.o(intermediate_reg_1[4370]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8739]),.i2(intermediate_reg_0[8738]),.o(intermediate_reg_1[4369])); 
fsm fsm_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8737]),.i2(intermediate_reg_0[8736]),.o(intermediate_reg_1[4368])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8735]),.i2(intermediate_reg_0[8734]),.o(intermediate_reg_1[4367]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8733]),.i2(intermediate_reg_0[8732]),.o(intermediate_reg_1[4366])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8731]),.i2(intermediate_reg_0[8730]),.o(intermediate_reg_1[4365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8729]),.i2(intermediate_reg_0[8728]),.o(intermediate_reg_1[4364]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8727]),.i2(intermediate_reg_0[8726]),.o(intermediate_reg_1[4363]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8725]),.i2(intermediate_reg_0[8724]),.o(intermediate_reg_1[4362]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8723]),.i2(intermediate_reg_0[8722]),.o(intermediate_reg_1[4361]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8721]),.i2(intermediate_reg_0[8720]),.o(intermediate_reg_1[4360])); 
fsm fsm_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8719]),.i2(intermediate_reg_0[8718]),.o(intermediate_reg_1[4359])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8717]),.i2(intermediate_reg_0[8716]),.o(intermediate_reg_1[4358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8715]),.i2(intermediate_reg_0[8714]),.o(intermediate_reg_1[4357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8713]),.i2(intermediate_reg_0[8712]),.o(intermediate_reg_1[4356]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8711]),.i2(intermediate_reg_0[8710]),.o(intermediate_reg_1[4355])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8709]),.i2(intermediate_reg_0[8708]),.o(intermediate_reg_1[4354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8707]),.i2(intermediate_reg_0[8706]),.o(intermediate_reg_1[4353]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8705]),.i2(intermediate_reg_0[8704]),.o(intermediate_reg_1[4352])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8703]),.i2(intermediate_reg_0[8702]),.o(intermediate_reg_1[4351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8701]),.i2(intermediate_reg_0[8700]),.o(intermediate_reg_1[4350]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8699]),.i2(intermediate_reg_0[8698]),.o(intermediate_reg_1[4349]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8697]),.i2(intermediate_reg_0[8696]),.o(intermediate_reg_1[4348]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8695]),.i2(intermediate_reg_0[8694]),.o(intermediate_reg_1[4347]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8693]),.i2(intermediate_reg_0[8692]),.o(intermediate_reg_1[4346])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8691]),.i2(intermediate_reg_0[8690]),.o(intermediate_reg_1[4345]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8689]),.i2(intermediate_reg_0[8688]),.o(intermediate_reg_1[4344])); 
fsm fsm_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8687]),.i2(intermediate_reg_0[8686]),.o(intermediate_reg_1[4343])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8685]),.i2(intermediate_reg_0[8684]),.o(intermediate_reg_1[4342]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8683]),.i2(intermediate_reg_0[8682]),.o(intermediate_reg_1[4341])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8681]),.i2(intermediate_reg_0[8680]),.o(intermediate_reg_1[4340])); 
mux_module mux_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8679]),.i2(intermediate_reg_0[8678]),.o(intermediate_reg_1[4339]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8677]),.i2(intermediate_reg_0[8676]),.o(intermediate_reg_1[4338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8675]),.i2(intermediate_reg_0[8674]),.o(intermediate_reg_1[4337]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8673]),.i2(intermediate_reg_0[8672]),.o(intermediate_reg_1[4336])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8671]),.i2(intermediate_reg_0[8670]),.o(intermediate_reg_1[4335])); 
mux_module mux_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8669]),.i2(intermediate_reg_0[8668]),.o(intermediate_reg_1[4334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8667]),.i2(intermediate_reg_0[8666]),.o(intermediate_reg_1[4333]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8665]),.i2(intermediate_reg_0[8664]),.o(intermediate_reg_1[4332])); 
mux_module mux_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8663]),.i2(intermediate_reg_0[8662]),.o(intermediate_reg_1[4331]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8661]),.i2(intermediate_reg_0[8660]),.o(intermediate_reg_1[4330])); 
fsm fsm_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8659]),.i2(intermediate_reg_0[8658]),.o(intermediate_reg_1[4329])); 
fsm fsm_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8657]),.i2(intermediate_reg_0[8656]),.o(intermediate_reg_1[4328])); 
mux_module mux_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8655]),.i2(intermediate_reg_0[8654]),.o(intermediate_reg_1[4327]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8653]),.i2(intermediate_reg_0[8652]),.o(intermediate_reg_1[4326]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8651]),.i2(intermediate_reg_0[8650]),.o(intermediate_reg_1[4325])); 
fsm fsm_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8649]),.i2(intermediate_reg_0[8648]),.o(intermediate_reg_1[4324])); 
fsm fsm_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8647]),.i2(intermediate_reg_0[8646]),.o(intermediate_reg_1[4323])); 
mux_module mux_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8645]),.i2(intermediate_reg_0[8644]),.o(intermediate_reg_1[4322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8643]),.i2(intermediate_reg_0[8642]),.o(intermediate_reg_1[4321]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8641]),.i2(intermediate_reg_0[8640]),.o(intermediate_reg_1[4320]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8639]),.i2(intermediate_reg_0[8638]),.o(intermediate_reg_1[4319])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8637]),.i2(intermediate_reg_0[8636]),.o(intermediate_reg_1[4318]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8635]),.i2(intermediate_reg_0[8634]),.o(intermediate_reg_1[4317])); 
fsm fsm_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8633]),.i2(intermediate_reg_0[8632]),.o(intermediate_reg_1[4316])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8631]),.i2(intermediate_reg_0[8630]),.o(intermediate_reg_1[4315]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8629]),.i2(intermediate_reg_0[8628]),.o(intermediate_reg_1[4314]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8627]),.i2(intermediate_reg_0[8626]),.o(intermediate_reg_1[4313])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8625]),.i2(intermediate_reg_0[8624]),.o(intermediate_reg_1[4312])); 
mux_module mux_module_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8623]),.i2(intermediate_reg_0[8622]),.o(intermediate_reg_1[4311]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8621]),.i2(intermediate_reg_0[8620]),.o(intermediate_reg_1[4310])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8619]),.i2(intermediate_reg_0[8618]),.o(intermediate_reg_1[4309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8617]),.i2(intermediate_reg_0[8616]),.o(intermediate_reg_1[4308]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8615]),.i2(intermediate_reg_0[8614]),.o(intermediate_reg_1[4307]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8613]),.i2(intermediate_reg_0[8612]),.o(intermediate_reg_1[4306])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8611]),.i2(intermediate_reg_0[8610]),.o(intermediate_reg_1[4305]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8609]),.i2(intermediate_reg_0[8608]),.o(intermediate_reg_1[4304])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8607]),.i2(intermediate_reg_0[8606]),.o(intermediate_reg_1[4303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8605]),.i2(intermediate_reg_0[8604]),.o(intermediate_reg_1[4302]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8603]),.i2(intermediate_reg_0[8602]),.o(intermediate_reg_1[4301])); 
fsm fsm_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8601]),.i2(intermediate_reg_0[8600]),.o(intermediate_reg_1[4300])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8599]),.i2(intermediate_reg_0[8598]),.o(intermediate_reg_1[4299]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8597]),.i2(intermediate_reg_0[8596]),.o(intermediate_reg_1[4298])); 
mux_module mux_module_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8595]),.i2(intermediate_reg_0[8594]),.o(intermediate_reg_1[4297]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8593]),.i2(intermediate_reg_0[8592]),.o(intermediate_reg_1[4296])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8591]),.i2(intermediate_reg_0[8590]),.o(intermediate_reg_1[4295]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8589]),.i2(intermediate_reg_0[8588]),.o(intermediate_reg_1[4294]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8587]),.i2(intermediate_reg_0[8586]),.o(intermediate_reg_1[4293]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8585]),.i2(intermediate_reg_0[8584]),.o(intermediate_reg_1[4292])); 
mux_module mux_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8583]),.i2(intermediate_reg_0[8582]),.o(intermediate_reg_1[4291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8581]),.i2(intermediate_reg_0[8580]),.o(intermediate_reg_1[4290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8579]),.i2(intermediate_reg_0[8578]),.o(intermediate_reg_1[4289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8577]),.i2(intermediate_reg_0[8576]),.o(intermediate_reg_1[4288]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8575]),.i2(intermediate_reg_0[8574]),.o(intermediate_reg_1[4287]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8573]),.i2(intermediate_reg_0[8572]),.o(intermediate_reg_1[4286])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8571]),.i2(intermediate_reg_0[8570]),.o(intermediate_reg_1[4285]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8569]),.i2(intermediate_reg_0[8568]),.o(intermediate_reg_1[4284])); 
fsm fsm_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8567]),.i2(intermediate_reg_0[8566]),.o(intermediate_reg_1[4283])); 
fsm fsm_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8565]),.i2(intermediate_reg_0[8564]),.o(intermediate_reg_1[4282])); 
fsm fsm_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8563]),.i2(intermediate_reg_0[8562]),.o(intermediate_reg_1[4281])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8561]),.i2(intermediate_reg_0[8560]),.o(intermediate_reg_1[4280])); 
fsm fsm_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8559]),.i2(intermediate_reg_0[8558]),.o(intermediate_reg_1[4279])); 
fsm fsm_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8557]),.i2(intermediate_reg_0[8556]),.o(intermediate_reg_1[4278])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8555]),.i2(intermediate_reg_0[8554]),.o(intermediate_reg_1[4277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8553]),.i2(intermediate_reg_0[8552]),.o(intermediate_reg_1[4276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8551]),.i2(intermediate_reg_0[8550]),.o(intermediate_reg_1[4275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8549]),.i2(intermediate_reg_0[8548]),.o(intermediate_reg_1[4274]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8547]),.i2(intermediate_reg_0[8546]),.o(intermediate_reg_1[4273])); 
mux_module mux_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8545]),.i2(intermediate_reg_0[8544]),.o(intermediate_reg_1[4272]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8543]),.i2(intermediate_reg_0[8542]),.o(intermediate_reg_1[4271])); 
mux_module mux_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8541]),.i2(intermediate_reg_0[8540]),.o(intermediate_reg_1[4270]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8539]),.i2(intermediate_reg_0[8538]),.o(intermediate_reg_1[4269])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8537]),.i2(intermediate_reg_0[8536]),.o(intermediate_reg_1[4268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8535]),.i2(intermediate_reg_0[8534]),.o(intermediate_reg_1[4267]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8533]),.i2(intermediate_reg_0[8532]),.o(intermediate_reg_1[4266]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8531]),.i2(intermediate_reg_0[8530]),.o(intermediate_reg_1[4265])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8529]),.i2(intermediate_reg_0[8528]),.o(intermediate_reg_1[4264]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8527]),.i2(intermediate_reg_0[8526]),.o(intermediate_reg_1[4263])); 
fsm fsm_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8525]),.i2(intermediate_reg_0[8524]),.o(intermediate_reg_1[4262])); 
mux_module mux_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8523]),.i2(intermediate_reg_0[8522]),.o(intermediate_reg_1[4261]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8521]),.i2(intermediate_reg_0[8520]),.o(intermediate_reg_1[4260])); 
fsm fsm_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8519]),.i2(intermediate_reg_0[8518]),.o(intermediate_reg_1[4259])); 
fsm fsm_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8517]),.i2(intermediate_reg_0[8516]),.o(intermediate_reg_1[4258])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8515]),.i2(intermediate_reg_0[8514]),.o(intermediate_reg_1[4257]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8513]),.i2(intermediate_reg_0[8512]),.o(intermediate_reg_1[4256])); 
fsm fsm_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8511]),.i2(intermediate_reg_0[8510]),.o(intermediate_reg_1[4255])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8509]),.i2(intermediate_reg_0[8508]),.o(intermediate_reg_1[4254])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8507]),.i2(intermediate_reg_0[8506]),.o(intermediate_reg_1[4253]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8505]),.i2(intermediate_reg_0[8504]),.o(intermediate_reg_1[4252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8503]),.i2(intermediate_reg_0[8502]),.o(intermediate_reg_1[4251]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8501]),.i2(intermediate_reg_0[8500]),.o(intermediate_reg_1[4250])); 
fsm fsm_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8499]),.i2(intermediate_reg_0[8498]),.o(intermediate_reg_1[4249])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8497]),.i2(intermediate_reg_0[8496]),.o(intermediate_reg_1[4248])); 
fsm fsm_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8495]),.i2(intermediate_reg_0[8494]),.o(intermediate_reg_1[4247])); 
mux_module mux_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8493]),.i2(intermediate_reg_0[8492]),.o(intermediate_reg_1[4246]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8491]),.i2(intermediate_reg_0[8490]),.o(intermediate_reg_1[4245])); 
mux_module mux_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8489]),.i2(intermediate_reg_0[8488]),.o(intermediate_reg_1[4244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8487]),.i2(intermediate_reg_0[8486]),.o(intermediate_reg_1[4243]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8485]),.i2(intermediate_reg_0[8484]),.o(intermediate_reg_1[4242])); 
mux_module mux_module_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8483]),.i2(intermediate_reg_0[8482]),.o(intermediate_reg_1[4241]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8481]),.i2(intermediate_reg_0[8480]),.o(intermediate_reg_1[4240])); 
fsm fsm_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8479]),.i2(intermediate_reg_0[8478]),.o(intermediate_reg_1[4239])); 
fsm fsm_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8477]),.i2(intermediate_reg_0[8476]),.o(intermediate_reg_1[4238])); 
fsm fsm_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8475]),.i2(intermediate_reg_0[8474]),.o(intermediate_reg_1[4237])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8473]),.i2(intermediate_reg_0[8472]),.o(intermediate_reg_1[4236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8471]),.i2(intermediate_reg_0[8470]),.o(intermediate_reg_1[4235]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8469]),.i2(intermediate_reg_0[8468]),.o(intermediate_reg_1[4234])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8467]),.i2(intermediate_reg_0[8466]),.o(intermediate_reg_1[4233]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8465]),.i2(intermediate_reg_0[8464]),.o(intermediate_reg_1[4232])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8463]),.i2(intermediate_reg_0[8462]),.o(intermediate_reg_1[4231]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8461]),.i2(intermediate_reg_0[8460]),.o(intermediate_reg_1[4230]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8459]),.i2(intermediate_reg_0[8458]),.o(intermediate_reg_1[4229])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8457]),.i2(intermediate_reg_0[8456]),.o(intermediate_reg_1[4228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8455]),.i2(intermediate_reg_0[8454]),.o(intermediate_reg_1[4227]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8453]),.i2(intermediate_reg_0[8452]),.o(intermediate_reg_1[4226])); 
fsm fsm_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8451]),.i2(intermediate_reg_0[8450]),.o(intermediate_reg_1[4225])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8449]),.i2(intermediate_reg_0[8448]),.o(intermediate_reg_1[4224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8447]),.i2(intermediate_reg_0[8446]),.o(intermediate_reg_1[4223]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8445]),.i2(intermediate_reg_0[8444]),.o(intermediate_reg_1[4222]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8443]),.i2(intermediate_reg_0[8442]),.o(intermediate_reg_1[4221]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8441]),.i2(intermediate_reg_0[8440]),.o(intermediate_reg_1[4220]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8439]),.i2(intermediate_reg_0[8438]),.o(intermediate_reg_1[4219])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8437]),.i2(intermediate_reg_0[8436]),.o(intermediate_reg_1[4218]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8435]),.i2(intermediate_reg_0[8434]),.o(intermediate_reg_1[4217])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8433]),.i2(intermediate_reg_0[8432]),.o(intermediate_reg_1[4216]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8431]),.i2(intermediate_reg_0[8430]),.o(intermediate_reg_1[4215])); 
mux_module mux_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8429]),.i2(intermediate_reg_0[8428]),.o(intermediate_reg_1[4214]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8427]),.i2(intermediate_reg_0[8426]),.o(intermediate_reg_1[4213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8425]),.i2(intermediate_reg_0[8424]),.o(intermediate_reg_1[4212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8423]),.i2(intermediate_reg_0[8422]),.o(intermediate_reg_1[4211]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8421]),.i2(intermediate_reg_0[8420]),.o(intermediate_reg_1[4210])); 
fsm fsm_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8419]),.i2(intermediate_reg_0[8418]),.o(intermediate_reg_1[4209])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8417]),.i2(intermediate_reg_0[8416]),.o(intermediate_reg_1[4208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8415]),.i2(intermediate_reg_0[8414]),.o(intermediate_reg_1[4207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8413]),.i2(intermediate_reg_0[8412]),.o(intermediate_reg_1[4206]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8411]),.i2(intermediate_reg_0[8410]),.o(intermediate_reg_1[4205])); 
mux_module mux_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8409]),.i2(intermediate_reg_0[8408]),.o(intermediate_reg_1[4204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8407]),.i2(intermediate_reg_0[8406]),.o(intermediate_reg_1[4203]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8405]),.i2(intermediate_reg_0[8404]),.o(intermediate_reg_1[4202])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8403]),.i2(intermediate_reg_0[8402]),.o(intermediate_reg_1[4201]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8401]),.i2(intermediate_reg_0[8400]),.o(intermediate_reg_1[4200])); 
mux_module mux_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8399]),.i2(intermediate_reg_0[8398]),.o(intermediate_reg_1[4199]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8397]),.i2(intermediate_reg_0[8396]),.o(intermediate_reg_1[4198]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8395]),.i2(intermediate_reg_0[8394]),.o(intermediate_reg_1[4197])); 
fsm fsm_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8393]),.i2(intermediate_reg_0[8392]),.o(intermediate_reg_1[4196])); 
fsm fsm_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8391]),.i2(intermediate_reg_0[8390]),.o(intermediate_reg_1[4195])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8389]),.i2(intermediate_reg_0[8388]),.o(intermediate_reg_1[4194]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8387]),.i2(intermediate_reg_0[8386]),.o(intermediate_reg_1[4193])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8385]),.i2(intermediate_reg_0[8384]),.o(intermediate_reg_1[4192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8383]),.i2(intermediate_reg_0[8382]),.o(intermediate_reg_1[4191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8381]),.i2(intermediate_reg_0[8380]),.o(intermediate_reg_1[4190]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8379]),.i2(intermediate_reg_0[8378]),.o(intermediate_reg_1[4189])); 
mux_module mux_module_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8377]),.i2(intermediate_reg_0[8376]),.o(intermediate_reg_1[4188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8375]),.i2(intermediate_reg_0[8374]),.o(intermediate_reg_1[4187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8373]),.i2(intermediate_reg_0[8372]),.o(intermediate_reg_1[4186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8371]),.i2(intermediate_reg_0[8370]),.o(intermediate_reg_1[4185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8369]),.i2(intermediate_reg_0[8368]),.o(intermediate_reg_1[4184]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8367]),.i2(intermediate_reg_0[8366]),.o(intermediate_reg_1[4183])); 
fsm fsm_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8365]),.i2(intermediate_reg_0[8364]),.o(intermediate_reg_1[4182])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8363]),.i2(intermediate_reg_0[8362]),.o(intermediate_reg_1[4181]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8361]),.i2(intermediate_reg_0[8360]),.o(intermediate_reg_1[4180])); 
fsm fsm_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8359]),.i2(intermediate_reg_0[8358]),.o(intermediate_reg_1[4179])); 
fsm fsm_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8357]),.i2(intermediate_reg_0[8356]),.o(intermediate_reg_1[4178])); 
fsm fsm_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8355]),.i2(intermediate_reg_0[8354]),.o(intermediate_reg_1[4177])); 
fsm fsm_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8353]),.i2(intermediate_reg_0[8352]),.o(intermediate_reg_1[4176])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8351]),.i2(intermediate_reg_0[8350]),.o(intermediate_reg_1[4175]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8349]),.i2(intermediate_reg_0[8348]),.o(intermediate_reg_1[4174])); 
fsm fsm_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8347]),.i2(intermediate_reg_0[8346]),.o(intermediate_reg_1[4173])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8345]),.i2(intermediate_reg_0[8344]),.o(intermediate_reg_1[4172])); 
fsm fsm_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8343]),.i2(intermediate_reg_0[8342]),.o(intermediate_reg_1[4171])); 
mux_module mux_module_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8341]),.i2(intermediate_reg_0[8340]),.o(intermediate_reg_1[4170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8339]),.i2(intermediate_reg_0[8338]),.o(intermediate_reg_1[4169]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8337]),.i2(intermediate_reg_0[8336]),.o(intermediate_reg_1[4168])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8335]),.i2(intermediate_reg_0[8334]),.o(intermediate_reg_1[4167]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8333]),.i2(intermediate_reg_0[8332]),.o(intermediate_reg_1[4166])); 
fsm fsm_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8331]),.i2(intermediate_reg_0[8330]),.o(intermediate_reg_1[4165])); 
fsm fsm_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8329]),.i2(intermediate_reg_0[8328]),.o(intermediate_reg_1[4164])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8327]),.i2(intermediate_reg_0[8326]),.o(intermediate_reg_1[4163])); 
fsm fsm_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8325]),.i2(intermediate_reg_0[8324]),.o(intermediate_reg_1[4162])); 
mux_module mux_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8323]),.i2(intermediate_reg_0[8322]),.o(intermediate_reg_1[4161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8321]),.i2(intermediate_reg_0[8320]),.o(intermediate_reg_1[4160]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8319]),.i2(intermediate_reg_0[8318]),.o(intermediate_reg_1[4159])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8317]),.i2(intermediate_reg_0[8316]),.o(intermediate_reg_1[4158])); 
fsm fsm_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8315]),.i2(intermediate_reg_0[8314]),.o(intermediate_reg_1[4157])); 
fsm fsm_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8313]),.i2(intermediate_reg_0[8312]),.o(intermediate_reg_1[4156])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8311]),.i2(intermediate_reg_0[8310]),.o(intermediate_reg_1[4155]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8309]),.i2(intermediate_reg_0[8308]),.o(intermediate_reg_1[4154]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8307]),.i2(intermediate_reg_0[8306]),.o(intermediate_reg_1[4153])); 
mux_module mux_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8305]),.i2(intermediate_reg_0[8304]),.o(intermediate_reg_1[4152]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8303]),.i2(intermediate_reg_0[8302]),.o(intermediate_reg_1[4151])); 
fsm fsm_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8301]),.i2(intermediate_reg_0[8300]),.o(intermediate_reg_1[4150])); 
mux_module mux_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8299]),.i2(intermediate_reg_0[8298]),.o(intermediate_reg_1[4149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8297]),.i2(intermediate_reg_0[8296]),.o(intermediate_reg_1[4148]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8295]),.i2(intermediate_reg_0[8294]),.o(intermediate_reg_1[4147])); 
mux_module mux_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8293]),.i2(intermediate_reg_0[8292]),.o(intermediate_reg_1[4146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8291]),.i2(intermediate_reg_0[8290]),.o(intermediate_reg_1[4145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8289]),.i2(intermediate_reg_0[8288]),.o(intermediate_reg_1[4144]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8287]),.i2(intermediate_reg_0[8286]),.o(intermediate_reg_1[4143])); 
fsm fsm_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8285]),.i2(intermediate_reg_0[8284]),.o(intermediate_reg_1[4142])); 
fsm fsm_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8283]),.i2(intermediate_reg_0[8282]),.o(intermediate_reg_1[4141])); 
fsm fsm_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8281]),.i2(intermediate_reg_0[8280]),.o(intermediate_reg_1[4140])); 
mux_module mux_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8279]),.i2(intermediate_reg_0[8278]),.o(intermediate_reg_1[4139]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8277]),.i2(intermediate_reg_0[8276]),.o(intermediate_reg_1[4138])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8275]),.i2(intermediate_reg_0[8274]),.o(intermediate_reg_1[4137]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8273]),.i2(intermediate_reg_0[8272]),.o(intermediate_reg_1[4136])); 
fsm fsm_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8271]),.i2(intermediate_reg_0[8270]),.o(intermediate_reg_1[4135])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8269]),.i2(intermediate_reg_0[8268]),.o(intermediate_reg_1[4134]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8267]),.i2(intermediate_reg_0[8266]),.o(intermediate_reg_1[4133])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8265]),.i2(intermediate_reg_0[8264]),.o(intermediate_reg_1[4132]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8263]),.i2(intermediate_reg_0[8262]),.o(intermediate_reg_1[4131])); 
fsm fsm_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8261]),.i2(intermediate_reg_0[8260]),.o(intermediate_reg_1[4130])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8259]),.i2(intermediate_reg_0[8258]),.o(intermediate_reg_1[4129])); 
fsm fsm_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8257]),.i2(intermediate_reg_0[8256]),.o(intermediate_reg_1[4128])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8255]),.i2(intermediate_reg_0[8254]),.o(intermediate_reg_1[4127]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8253]),.i2(intermediate_reg_0[8252]),.o(intermediate_reg_1[4126])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8251]),.i2(intermediate_reg_0[8250]),.o(intermediate_reg_1[4125]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8249]),.i2(intermediate_reg_0[8248]),.o(intermediate_reg_1[4124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8247]),.i2(intermediate_reg_0[8246]),.o(intermediate_reg_1[4123]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8245]),.i2(intermediate_reg_0[8244]),.o(intermediate_reg_1[4122]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8243]),.i2(intermediate_reg_0[8242]),.o(intermediate_reg_1[4121])); 
mux_module mux_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8241]),.i2(intermediate_reg_0[8240]),.o(intermediate_reg_1[4120]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8239]),.i2(intermediate_reg_0[8238]),.o(intermediate_reg_1[4119])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8237]),.i2(intermediate_reg_0[8236]),.o(intermediate_reg_1[4118])); 
fsm fsm_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8235]),.i2(intermediate_reg_0[8234]),.o(intermediate_reg_1[4117])); 
fsm fsm_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8233]),.i2(intermediate_reg_0[8232]),.o(intermediate_reg_1[4116])); 
mux_module mux_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8231]),.i2(intermediate_reg_0[8230]),.o(intermediate_reg_1[4115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8229]),.i2(intermediate_reg_0[8228]),.o(intermediate_reg_1[4114])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8227]),.i2(intermediate_reg_0[8226]),.o(intermediate_reg_1[4113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8225]),.i2(intermediate_reg_0[8224]),.o(intermediate_reg_1[4112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8223]),.i2(intermediate_reg_0[8222]),.o(intermediate_reg_1[4111]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8221]),.i2(intermediate_reg_0[8220]),.o(intermediate_reg_1[4110]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8219]),.i2(intermediate_reg_0[8218]),.o(intermediate_reg_1[4109])); 
fsm fsm_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8217]),.i2(intermediate_reg_0[8216]),.o(intermediate_reg_1[4108])); 
fsm fsm_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8215]),.i2(intermediate_reg_0[8214]),.o(intermediate_reg_1[4107])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8213]),.i2(intermediate_reg_0[8212]),.o(intermediate_reg_1[4106]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8211]),.i2(intermediate_reg_0[8210]),.o(intermediate_reg_1[4105])); 
fsm fsm_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8209]),.i2(intermediate_reg_0[8208]),.o(intermediate_reg_1[4104])); 
mux_module mux_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8207]),.i2(intermediate_reg_0[8206]),.o(intermediate_reg_1[4103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8205]),.i2(intermediate_reg_0[8204]),.o(intermediate_reg_1[4102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8203]),.i2(intermediate_reg_0[8202]),.o(intermediate_reg_1[4101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8201]),.i2(intermediate_reg_0[8200]),.o(intermediate_reg_1[4100]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8199]),.i2(intermediate_reg_0[8198]),.o(intermediate_reg_1[4099])); 
fsm fsm_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8197]),.i2(intermediate_reg_0[8196]),.o(intermediate_reg_1[4098])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8195]),.i2(intermediate_reg_0[8194]),.o(intermediate_reg_1[4097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8193]),.i2(intermediate_reg_0[8192]),.o(intermediate_reg_1[4096]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8191]),.i2(intermediate_reg_0[8190]),.o(intermediate_reg_1[4095])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8189]),.i2(intermediate_reg_0[8188]),.o(intermediate_reg_1[4094]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8187]),.i2(intermediate_reg_0[8186]),.o(intermediate_reg_1[4093])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8185]),.i2(intermediate_reg_0[8184]),.o(intermediate_reg_1[4092]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8183]),.i2(intermediate_reg_0[8182]),.o(intermediate_reg_1[4091])); 
mux_module mux_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8181]),.i2(intermediate_reg_0[8180]),.o(intermediate_reg_1[4090]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8179]),.i2(intermediate_reg_0[8178]),.o(intermediate_reg_1[4089])); 
fsm fsm_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8177]),.i2(intermediate_reg_0[8176]),.o(intermediate_reg_1[4088])); 
fsm fsm_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8175]),.i2(intermediate_reg_0[8174]),.o(intermediate_reg_1[4087])); 
fsm fsm_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8173]),.i2(intermediate_reg_0[8172]),.o(intermediate_reg_1[4086])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8171]),.i2(intermediate_reg_0[8170]),.o(intermediate_reg_1[4085]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8169]),.i2(intermediate_reg_0[8168]),.o(intermediate_reg_1[4084]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8167]),.i2(intermediate_reg_0[8166]),.o(intermediate_reg_1[4083])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8165]),.i2(intermediate_reg_0[8164]),.o(intermediate_reg_1[4082])); 
fsm fsm_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8163]),.i2(intermediate_reg_0[8162]),.o(intermediate_reg_1[4081])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8161]),.i2(intermediate_reg_0[8160]),.o(intermediate_reg_1[4080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8159]),.i2(intermediate_reg_0[8158]),.o(intermediate_reg_1[4079]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8157]),.i2(intermediate_reg_0[8156]),.o(intermediate_reg_1[4078])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8155]),.i2(intermediate_reg_0[8154]),.o(intermediate_reg_1[4077])); 
fsm fsm_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8153]),.i2(intermediate_reg_0[8152]),.o(intermediate_reg_1[4076])); 
fsm fsm_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8151]),.i2(intermediate_reg_0[8150]),.o(intermediate_reg_1[4075])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8149]),.i2(intermediate_reg_0[8148]),.o(intermediate_reg_1[4074]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8147]),.i2(intermediate_reg_0[8146]),.o(intermediate_reg_1[4073])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8145]),.i2(intermediate_reg_0[8144]),.o(intermediate_reg_1[4072]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8143]),.i2(intermediate_reg_0[8142]),.o(intermediate_reg_1[4071]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8141]),.i2(intermediate_reg_0[8140]),.o(intermediate_reg_1[4070]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8139]),.i2(intermediate_reg_0[8138]),.o(intermediate_reg_1[4069])); 
fsm fsm_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8137]),.i2(intermediate_reg_0[8136]),.o(intermediate_reg_1[4068])); 
fsm fsm_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8135]),.i2(intermediate_reg_0[8134]),.o(intermediate_reg_1[4067])); 
fsm fsm_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8133]),.i2(intermediate_reg_0[8132]),.o(intermediate_reg_1[4066])); 
fsm fsm_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8131]),.i2(intermediate_reg_0[8130]),.o(intermediate_reg_1[4065])); 
fsm fsm_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8129]),.i2(intermediate_reg_0[8128]),.o(intermediate_reg_1[4064])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8127]),.i2(intermediate_reg_0[8126]),.o(intermediate_reg_1[4063])); 
mux_module mux_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8125]),.i2(intermediate_reg_0[8124]),.o(intermediate_reg_1[4062]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8123]),.i2(intermediate_reg_0[8122]),.o(intermediate_reg_1[4061])); 
mux_module mux_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8121]),.i2(intermediate_reg_0[8120]),.o(intermediate_reg_1[4060]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8119]),.i2(intermediate_reg_0[8118]),.o(intermediate_reg_1[4059])); 
fsm fsm_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8117]),.i2(intermediate_reg_0[8116]),.o(intermediate_reg_1[4058])); 
fsm fsm_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8115]),.i2(intermediate_reg_0[8114]),.o(intermediate_reg_1[4057])); 
mux_module mux_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8113]),.i2(intermediate_reg_0[8112]),.o(intermediate_reg_1[4056]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8111]),.i2(intermediate_reg_0[8110]),.o(intermediate_reg_1[4055])); 
fsm fsm_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8109]),.i2(intermediate_reg_0[8108]),.o(intermediate_reg_1[4054])); 
fsm fsm_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8107]),.i2(intermediate_reg_0[8106]),.o(intermediate_reg_1[4053])); 
mux_module mux_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8105]),.i2(intermediate_reg_0[8104]),.o(intermediate_reg_1[4052]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8103]),.i2(intermediate_reg_0[8102]),.o(intermediate_reg_1[4051])); 
fsm fsm_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8101]),.i2(intermediate_reg_0[8100]),.o(intermediate_reg_1[4050])); 
fsm fsm_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8099]),.i2(intermediate_reg_0[8098]),.o(intermediate_reg_1[4049])); 
mux_module mux_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8097]),.i2(intermediate_reg_0[8096]),.o(intermediate_reg_1[4048]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8095]),.i2(intermediate_reg_0[8094]),.o(intermediate_reg_1[4047])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8093]),.i2(intermediate_reg_0[8092]),.o(intermediate_reg_1[4046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8091]),.i2(intermediate_reg_0[8090]),.o(intermediate_reg_1[4045]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8089]),.i2(intermediate_reg_0[8088]),.o(intermediate_reg_1[4044])); 
fsm fsm_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8087]),.i2(intermediate_reg_0[8086]),.o(intermediate_reg_1[4043])); 
fsm fsm_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8085]),.i2(intermediate_reg_0[8084]),.o(intermediate_reg_1[4042])); 
fsm fsm_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8083]),.i2(intermediate_reg_0[8082]),.o(intermediate_reg_1[4041])); 
fsm fsm_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8081]),.i2(intermediate_reg_0[8080]),.o(intermediate_reg_1[4040])); 
fsm fsm_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8079]),.i2(intermediate_reg_0[8078]),.o(intermediate_reg_1[4039])); 
fsm fsm_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8077]),.i2(intermediate_reg_0[8076]),.o(intermediate_reg_1[4038])); 
mux_module mux_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8075]),.i2(intermediate_reg_0[8074]),.o(intermediate_reg_1[4037]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8073]),.i2(intermediate_reg_0[8072]),.o(intermediate_reg_1[4036]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8071]),.i2(intermediate_reg_0[8070]),.o(intermediate_reg_1[4035])); 
mux_module mux_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8069]),.i2(intermediate_reg_0[8068]),.o(intermediate_reg_1[4034]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8067]),.i2(intermediate_reg_0[8066]),.o(intermediate_reg_1[4033]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8065]),.i2(intermediate_reg_0[8064]),.o(intermediate_reg_1[4032]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8063]),.i2(intermediate_reg_0[8062]),.o(intermediate_reg_1[4031])); 
fsm fsm_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8061]),.i2(intermediate_reg_0[8060]),.o(intermediate_reg_1[4030])); 
mux_module mux_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8059]),.i2(intermediate_reg_0[8058]),.o(intermediate_reg_1[4029]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8057]),.i2(intermediate_reg_0[8056]),.o(intermediate_reg_1[4028])); 
mux_module mux_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8055]),.i2(intermediate_reg_0[8054]),.o(intermediate_reg_1[4027]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8053]),.i2(intermediate_reg_0[8052]),.o(intermediate_reg_1[4026])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8051]),.i2(intermediate_reg_0[8050]),.o(intermediate_reg_1[4025])); 
fsm fsm_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8049]),.i2(intermediate_reg_0[8048]),.o(intermediate_reg_1[4024])); 
fsm fsm_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8047]),.i2(intermediate_reg_0[8046]),.o(intermediate_reg_1[4023])); 
mux_module mux_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8045]),.i2(intermediate_reg_0[8044]),.o(intermediate_reg_1[4022]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8043]),.i2(intermediate_reg_0[8042]),.o(intermediate_reg_1[4021])); 
fsm fsm_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8041]),.i2(intermediate_reg_0[8040]),.o(intermediate_reg_1[4020])); 
fsm fsm_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8039]),.i2(intermediate_reg_0[8038]),.o(intermediate_reg_1[4019])); 
fsm fsm_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8037]),.i2(intermediate_reg_0[8036]),.o(intermediate_reg_1[4018])); 
mux_module mux_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8035]),.i2(intermediate_reg_0[8034]),.o(intermediate_reg_1[4017]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8033]),.i2(intermediate_reg_0[8032]),.o(intermediate_reg_1[4016]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8031]),.i2(intermediate_reg_0[8030]),.o(intermediate_reg_1[4015]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8029]),.i2(intermediate_reg_0[8028]),.o(intermediate_reg_1[4014]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8027]),.i2(intermediate_reg_0[8026]),.o(intermediate_reg_1[4013])); 
fsm fsm_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8025]),.i2(intermediate_reg_0[8024]),.o(intermediate_reg_1[4012])); 
mux_module mux_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8023]),.i2(intermediate_reg_0[8022]),.o(intermediate_reg_1[4011]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8021]),.i2(intermediate_reg_0[8020]),.o(intermediate_reg_1[4010])); 
mux_module mux_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8019]),.i2(intermediate_reg_0[8018]),.o(intermediate_reg_1[4009]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8017]),.i2(intermediate_reg_0[8016]),.o(intermediate_reg_1[4008]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8015]),.i2(intermediate_reg_0[8014]),.o(intermediate_reg_1[4007]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8013]),.i2(intermediate_reg_0[8012]),.o(intermediate_reg_1[4006])); 
fsm fsm_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8011]),.i2(intermediate_reg_0[8010]),.o(intermediate_reg_1[4005])); 
fsm fsm_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8009]),.i2(intermediate_reg_0[8008]),.o(intermediate_reg_1[4004])); 
mux_module mux_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8007]),.i2(intermediate_reg_0[8006]),.o(intermediate_reg_1[4003]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8005]),.i2(intermediate_reg_0[8004]),.o(intermediate_reg_1[4002]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8003]),.i2(intermediate_reg_0[8002]),.o(intermediate_reg_1[4001])); 
fsm fsm_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[8001]),.i2(intermediate_reg_0[8000]),.o(intermediate_reg_1[4000])); 
fsm fsm_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7999]),.i2(intermediate_reg_0[7998]),.o(intermediate_reg_1[3999])); 
mux_module mux_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7997]),.i2(intermediate_reg_0[7996]),.o(intermediate_reg_1[3998]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7995]),.i2(intermediate_reg_0[7994]),.o(intermediate_reg_1[3997])); 
fsm fsm_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7993]),.i2(intermediate_reg_0[7992]),.o(intermediate_reg_1[3996])); 
mux_module mux_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7991]),.i2(intermediate_reg_0[7990]),.o(intermediate_reg_1[3995]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7989]),.i2(intermediate_reg_0[7988]),.o(intermediate_reg_1[3994]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7987]),.i2(intermediate_reg_0[7986]),.o(intermediate_reg_1[3993])); 
fsm fsm_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7985]),.i2(intermediate_reg_0[7984]),.o(intermediate_reg_1[3992])); 
mux_module mux_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7983]),.i2(intermediate_reg_0[7982]),.o(intermediate_reg_1[3991]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7981]),.i2(intermediate_reg_0[7980]),.o(intermediate_reg_1[3990])); 
fsm fsm_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7979]),.i2(intermediate_reg_0[7978]),.o(intermediate_reg_1[3989])); 
fsm fsm_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7977]),.i2(intermediate_reg_0[7976]),.o(intermediate_reg_1[3988])); 
mux_module mux_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7975]),.i2(intermediate_reg_0[7974]),.o(intermediate_reg_1[3987]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7973]),.i2(intermediate_reg_0[7972]),.o(intermediate_reg_1[3986]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7971]),.i2(intermediate_reg_0[7970]),.o(intermediate_reg_1[3985])); 
fsm fsm_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7969]),.i2(intermediate_reg_0[7968]),.o(intermediate_reg_1[3984])); 
mux_module mux_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7967]),.i2(intermediate_reg_0[7966]),.o(intermediate_reg_1[3983]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7965]),.i2(intermediate_reg_0[7964]),.o(intermediate_reg_1[3982])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7963]),.i2(intermediate_reg_0[7962]),.o(intermediate_reg_1[3981]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7961]),.i2(intermediate_reg_0[7960]),.o(intermediate_reg_1[3980])); 
fsm fsm_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7959]),.i2(intermediate_reg_0[7958]),.o(intermediate_reg_1[3979])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7957]),.i2(intermediate_reg_0[7956]),.o(intermediate_reg_1[3978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7955]),.i2(intermediate_reg_0[7954]),.o(intermediate_reg_1[3977]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7953]),.i2(intermediate_reg_0[7952]),.o(intermediate_reg_1[3976])); 
mux_module mux_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7951]),.i2(intermediate_reg_0[7950]),.o(intermediate_reg_1[3975]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7949]),.i2(intermediate_reg_0[7948]),.o(intermediate_reg_1[3974])); 
fsm fsm_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7947]),.i2(intermediate_reg_0[7946]),.o(intermediate_reg_1[3973])); 
fsm fsm_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7945]),.i2(intermediate_reg_0[7944]),.o(intermediate_reg_1[3972])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7943]),.i2(intermediate_reg_0[7942]),.o(intermediate_reg_1[3971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7941]),.i2(intermediate_reg_0[7940]),.o(intermediate_reg_1[3970]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7939]),.i2(intermediate_reg_0[7938]),.o(intermediate_reg_1[3969])); 
fsm fsm_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7937]),.i2(intermediate_reg_0[7936]),.o(intermediate_reg_1[3968])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7935]),.i2(intermediate_reg_0[7934]),.o(intermediate_reg_1[3967]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7933]),.i2(intermediate_reg_0[7932]),.o(intermediate_reg_1[3966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7931]),.i2(intermediate_reg_0[7930]),.o(intermediate_reg_1[3965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7929]),.i2(intermediate_reg_0[7928]),.o(intermediate_reg_1[3964]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7927]),.i2(intermediate_reg_0[7926]),.o(intermediate_reg_1[3963])); 
fsm fsm_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7925]),.i2(intermediate_reg_0[7924]),.o(intermediate_reg_1[3962])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7923]),.i2(intermediate_reg_0[7922]),.o(intermediate_reg_1[3961]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7921]),.i2(intermediate_reg_0[7920]),.o(intermediate_reg_1[3960])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7919]),.i2(intermediate_reg_0[7918]),.o(intermediate_reg_1[3959]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7917]),.i2(intermediate_reg_0[7916]),.o(intermediate_reg_1[3958]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7915]),.i2(intermediate_reg_0[7914]),.o(intermediate_reg_1[3957]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7913]),.i2(intermediate_reg_0[7912]),.o(intermediate_reg_1[3956])); 
mux_module mux_module_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7911]),.i2(intermediate_reg_0[7910]),.o(intermediate_reg_1[3955]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7909]),.i2(intermediate_reg_0[7908]),.o(intermediate_reg_1[3954]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7907]),.i2(intermediate_reg_0[7906]),.o(intermediate_reg_1[3953]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7905]),.i2(intermediate_reg_0[7904]),.o(intermediate_reg_1[3952]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7903]),.i2(intermediate_reg_0[7902]),.o(intermediate_reg_1[3951])); 
fsm fsm_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7901]),.i2(intermediate_reg_0[7900]),.o(intermediate_reg_1[3950])); 
mux_module mux_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7899]),.i2(intermediate_reg_0[7898]),.o(intermediate_reg_1[3949]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7897]),.i2(intermediate_reg_0[7896]),.o(intermediate_reg_1[3948])); 
fsm fsm_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7895]),.i2(intermediate_reg_0[7894]),.o(intermediate_reg_1[3947])); 
fsm fsm_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7893]),.i2(intermediate_reg_0[7892]),.o(intermediate_reg_1[3946])); 
fsm fsm_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7891]),.i2(intermediate_reg_0[7890]),.o(intermediate_reg_1[3945])); 
mux_module mux_module_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7889]),.i2(intermediate_reg_0[7888]),.o(intermediate_reg_1[3944]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7887]),.i2(intermediate_reg_0[7886]),.o(intermediate_reg_1[3943])); 
fsm fsm_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7885]),.i2(intermediate_reg_0[7884]),.o(intermediate_reg_1[3942])); 
fsm fsm_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7883]),.i2(intermediate_reg_0[7882]),.o(intermediate_reg_1[3941])); 
mux_module mux_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7881]),.i2(intermediate_reg_0[7880]),.o(intermediate_reg_1[3940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7879]),.i2(intermediate_reg_0[7878]),.o(intermediate_reg_1[3939]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7877]),.i2(intermediate_reg_0[7876]),.o(intermediate_reg_1[3938]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7875]),.i2(intermediate_reg_0[7874]),.o(intermediate_reg_1[3937]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7873]),.i2(intermediate_reg_0[7872]),.o(intermediate_reg_1[3936]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7871]),.i2(intermediate_reg_0[7870]),.o(intermediate_reg_1[3935])); 
fsm fsm_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7869]),.i2(intermediate_reg_0[7868]),.o(intermediate_reg_1[3934])); 
fsm fsm_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7867]),.i2(intermediate_reg_0[7866]),.o(intermediate_reg_1[3933])); 
fsm fsm_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7865]),.i2(intermediate_reg_0[7864]),.o(intermediate_reg_1[3932])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7863]),.i2(intermediate_reg_0[7862]),.o(intermediate_reg_1[3931]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7861]),.i2(intermediate_reg_0[7860]),.o(intermediate_reg_1[3930])); 
fsm fsm_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7859]),.i2(intermediate_reg_0[7858]),.o(intermediate_reg_1[3929])); 
mux_module mux_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7857]),.i2(intermediate_reg_0[7856]),.o(intermediate_reg_1[3928]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7855]),.i2(intermediate_reg_0[7854]),.o(intermediate_reg_1[3927])); 
mux_module mux_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7853]),.i2(intermediate_reg_0[7852]),.o(intermediate_reg_1[3926]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7851]),.i2(intermediate_reg_0[7850]),.o(intermediate_reg_1[3925])); 
fsm fsm_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7849]),.i2(intermediate_reg_0[7848]),.o(intermediate_reg_1[3924])); 
mux_module mux_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7847]),.i2(intermediate_reg_0[7846]),.o(intermediate_reg_1[3923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7845]),.i2(intermediate_reg_0[7844]),.o(intermediate_reg_1[3922]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7843]),.i2(intermediate_reg_0[7842]),.o(intermediate_reg_1[3921])); 
fsm fsm_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7841]),.i2(intermediate_reg_0[7840]),.o(intermediate_reg_1[3920])); 
fsm fsm_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7839]),.i2(intermediate_reg_0[7838]),.o(intermediate_reg_1[3919])); 
mux_module mux_module_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7837]),.i2(intermediate_reg_0[7836]),.o(intermediate_reg_1[3918]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7835]),.i2(intermediate_reg_0[7834]),.o(intermediate_reg_1[3917]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7833]),.i2(intermediate_reg_0[7832]),.o(intermediate_reg_1[3916])); 
mux_module mux_module_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7831]),.i2(intermediate_reg_0[7830]),.o(intermediate_reg_1[3915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7829]),.i2(intermediate_reg_0[7828]),.o(intermediate_reg_1[3914]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7827]),.i2(intermediate_reg_0[7826]),.o(intermediate_reg_1[3913])); 
fsm fsm_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7825]),.i2(intermediate_reg_0[7824]),.o(intermediate_reg_1[3912])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7823]),.i2(intermediate_reg_0[7822]),.o(intermediate_reg_1[3911]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7821]),.i2(intermediate_reg_0[7820]),.o(intermediate_reg_1[3910])); 
fsm fsm_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7819]),.i2(intermediate_reg_0[7818]),.o(intermediate_reg_1[3909])); 
fsm fsm_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7817]),.i2(intermediate_reg_0[7816]),.o(intermediate_reg_1[3908])); 
fsm fsm_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7815]),.i2(intermediate_reg_0[7814]),.o(intermediate_reg_1[3907])); 
fsm fsm_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7813]),.i2(intermediate_reg_0[7812]),.o(intermediate_reg_1[3906])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7811]),.i2(intermediate_reg_0[7810]),.o(intermediate_reg_1[3905]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7809]),.i2(intermediate_reg_0[7808]),.o(intermediate_reg_1[3904])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7807]),.i2(intermediate_reg_0[7806]),.o(intermediate_reg_1[3903]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7805]),.i2(intermediate_reg_0[7804]),.o(intermediate_reg_1[3902]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7803]),.i2(intermediate_reg_0[7802]),.o(intermediate_reg_1[3901]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7801]),.i2(intermediate_reg_0[7800]),.o(intermediate_reg_1[3900]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7799]),.i2(intermediate_reg_0[7798]),.o(intermediate_reg_1[3899])); 
fsm fsm_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7797]),.i2(intermediate_reg_0[7796]),.o(intermediate_reg_1[3898])); 
fsm fsm_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7795]),.i2(intermediate_reg_0[7794]),.o(intermediate_reg_1[3897])); 
fsm fsm_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7793]),.i2(intermediate_reg_0[7792]),.o(intermediate_reg_1[3896])); 
mux_module mux_module_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7791]),.i2(intermediate_reg_0[7790]),.o(intermediate_reg_1[3895]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7789]),.i2(intermediate_reg_0[7788]),.o(intermediate_reg_1[3894])); 
mux_module mux_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7787]),.i2(intermediate_reg_0[7786]),.o(intermediate_reg_1[3893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7785]),.i2(intermediate_reg_0[7784]),.o(intermediate_reg_1[3892]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7783]),.i2(intermediate_reg_0[7782]),.o(intermediate_reg_1[3891])); 
fsm fsm_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7781]),.i2(intermediate_reg_0[7780]),.o(intermediate_reg_1[3890])); 
mux_module mux_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7779]),.i2(intermediate_reg_0[7778]),.o(intermediate_reg_1[3889]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7777]),.i2(intermediate_reg_0[7776]),.o(intermediate_reg_1[3888])); 
mux_module mux_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7775]),.i2(intermediate_reg_0[7774]),.o(intermediate_reg_1[3887]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7773]),.i2(intermediate_reg_0[7772]),.o(intermediate_reg_1[3886])); 
mux_module mux_module_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7771]),.i2(intermediate_reg_0[7770]),.o(intermediate_reg_1[3885]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7769]),.i2(intermediate_reg_0[7768]),.o(intermediate_reg_1[3884])); 
mux_module mux_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7767]),.i2(intermediate_reg_0[7766]),.o(intermediate_reg_1[3883]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7765]),.i2(intermediate_reg_0[7764]),.o(intermediate_reg_1[3882])); 
mux_module mux_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7763]),.i2(intermediate_reg_0[7762]),.o(intermediate_reg_1[3881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7761]),.i2(intermediate_reg_0[7760]),.o(intermediate_reg_1[3880]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7759]),.i2(intermediate_reg_0[7758]),.o(intermediate_reg_1[3879])); 
mux_module mux_module_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7757]),.i2(intermediate_reg_0[7756]),.o(intermediate_reg_1[3878]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7755]),.i2(intermediate_reg_0[7754]),.o(intermediate_reg_1[3877]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7753]),.i2(intermediate_reg_0[7752]),.o(intermediate_reg_1[3876])); 
mux_module mux_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7751]),.i2(intermediate_reg_0[7750]),.o(intermediate_reg_1[3875]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7749]),.i2(intermediate_reg_0[7748]),.o(intermediate_reg_1[3874]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7747]),.i2(intermediate_reg_0[7746]),.o(intermediate_reg_1[3873]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7745]),.i2(intermediate_reg_0[7744]),.o(intermediate_reg_1[3872])); 
mux_module mux_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7743]),.i2(intermediate_reg_0[7742]),.o(intermediate_reg_1[3871]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7741]),.i2(intermediate_reg_0[7740]),.o(intermediate_reg_1[3870]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7739]),.i2(intermediate_reg_0[7738]),.o(intermediate_reg_1[3869])); 
fsm fsm_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7737]),.i2(intermediate_reg_0[7736]),.o(intermediate_reg_1[3868])); 
fsm fsm_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7735]),.i2(intermediate_reg_0[7734]),.o(intermediate_reg_1[3867])); 
mux_module mux_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7733]),.i2(intermediate_reg_0[7732]),.o(intermediate_reg_1[3866]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7731]),.i2(intermediate_reg_0[7730]),.o(intermediate_reg_1[3865])); 
mux_module mux_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7729]),.i2(intermediate_reg_0[7728]),.o(intermediate_reg_1[3864]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7727]),.i2(intermediate_reg_0[7726]),.o(intermediate_reg_1[3863])); 
mux_module mux_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7725]),.i2(intermediate_reg_0[7724]),.o(intermediate_reg_1[3862]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7723]),.i2(intermediate_reg_0[7722]),.o(intermediate_reg_1[3861]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7721]),.i2(intermediate_reg_0[7720]),.o(intermediate_reg_1[3860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7719]),.i2(intermediate_reg_0[7718]),.o(intermediate_reg_1[3859]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7717]),.i2(intermediate_reg_0[7716]),.o(intermediate_reg_1[3858]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7715]),.i2(intermediate_reg_0[7714]),.o(intermediate_reg_1[3857]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7713]),.i2(intermediate_reg_0[7712]),.o(intermediate_reg_1[3856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7711]),.i2(intermediate_reg_0[7710]),.o(intermediate_reg_1[3855]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7709]),.i2(intermediate_reg_0[7708]),.o(intermediate_reg_1[3854])); 
fsm fsm_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7707]),.i2(intermediate_reg_0[7706]),.o(intermediate_reg_1[3853])); 
fsm fsm_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7705]),.i2(intermediate_reg_0[7704]),.o(intermediate_reg_1[3852])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7703]),.i2(intermediate_reg_0[7702]),.o(intermediate_reg_1[3851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7701]),.i2(intermediate_reg_0[7700]),.o(intermediate_reg_1[3850]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7699]),.i2(intermediate_reg_0[7698]),.o(intermediate_reg_1[3849]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7697]),.i2(intermediate_reg_0[7696]),.o(intermediate_reg_1[3848])); 
mux_module mux_module_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7695]),.i2(intermediate_reg_0[7694]),.o(intermediate_reg_1[3847]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7693]),.i2(intermediate_reg_0[7692]),.o(intermediate_reg_1[3846])); 
fsm fsm_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7691]),.i2(intermediate_reg_0[7690]),.o(intermediate_reg_1[3845])); 
mux_module mux_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7689]),.i2(intermediate_reg_0[7688]),.o(intermediate_reg_1[3844]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7687]),.i2(intermediate_reg_0[7686]),.o(intermediate_reg_1[3843])); 
fsm fsm_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7685]),.i2(intermediate_reg_0[7684]),.o(intermediate_reg_1[3842])); 
mux_module mux_module_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7683]),.i2(intermediate_reg_0[7682]),.o(intermediate_reg_1[3841]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7681]),.i2(intermediate_reg_0[7680]),.o(intermediate_reg_1[3840])); 
mux_module mux_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7679]),.i2(intermediate_reg_0[7678]),.o(intermediate_reg_1[3839]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7677]),.i2(intermediate_reg_0[7676]),.o(intermediate_reg_1[3838]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7675]),.i2(intermediate_reg_0[7674]),.o(intermediate_reg_1[3837]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7673]),.i2(intermediate_reg_0[7672]),.o(intermediate_reg_1[3836]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7671]),.i2(intermediate_reg_0[7670]),.o(intermediate_reg_1[3835])); 
mux_module mux_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7669]),.i2(intermediate_reg_0[7668]),.o(intermediate_reg_1[3834]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7667]),.i2(intermediate_reg_0[7666]),.o(intermediate_reg_1[3833])); 
fsm fsm_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7665]),.i2(intermediate_reg_0[7664]),.o(intermediate_reg_1[3832])); 
fsm fsm_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7663]),.i2(intermediate_reg_0[7662]),.o(intermediate_reg_1[3831])); 
fsm fsm_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7661]),.i2(intermediate_reg_0[7660]),.o(intermediate_reg_1[3830])); 
mux_module mux_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7659]),.i2(intermediate_reg_0[7658]),.o(intermediate_reg_1[3829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7657]),.i2(intermediate_reg_0[7656]),.o(intermediate_reg_1[3828]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7655]),.i2(intermediate_reg_0[7654]),.o(intermediate_reg_1[3827])); 
mux_module mux_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7653]),.i2(intermediate_reg_0[7652]),.o(intermediate_reg_1[3826]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7651]),.i2(intermediate_reg_0[7650]),.o(intermediate_reg_1[3825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7649]),.i2(intermediate_reg_0[7648]),.o(intermediate_reg_1[3824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7647]),.i2(intermediate_reg_0[7646]),.o(intermediate_reg_1[3823]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7645]),.i2(intermediate_reg_0[7644]),.o(intermediate_reg_1[3822])); 
mux_module mux_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7643]),.i2(intermediate_reg_0[7642]),.o(intermediate_reg_1[3821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7641]),.i2(intermediate_reg_0[7640]),.o(intermediate_reg_1[3820]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7639]),.i2(intermediate_reg_0[7638]),.o(intermediate_reg_1[3819]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7637]),.i2(intermediate_reg_0[7636]),.o(intermediate_reg_1[3818])); 
fsm fsm_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7635]),.i2(intermediate_reg_0[7634]),.o(intermediate_reg_1[3817])); 
fsm fsm_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7633]),.i2(intermediate_reg_0[7632]),.o(intermediate_reg_1[3816])); 
mux_module mux_module_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7631]),.i2(intermediate_reg_0[7630]),.o(intermediate_reg_1[3815]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7629]),.i2(intermediate_reg_0[7628]),.o(intermediate_reg_1[3814])); 
mux_module mux_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7627]),.i2(intermediate_reg_0[7626]),.o(intermediate_reg_1[3813]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7625]),.i2(intermediate_reg_0[7624]),.o(intermediate_reg_1[3812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7623]),.i2(intermediate_reg_0[7622]),.o(intermediate_reg_1[3811]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7621]),.i2(intermediate_reg_0[7620]),.o(intermediate_reg_1[3810])); 
fsm fsm_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7619]),.i2(intermediate_reg_0[7618]),.o(intermediate_reg_1[3809])); 
mux_module mux_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7617]),.i2(intermediate_reg_0[7616]),.o(intermediate_reg_1[3808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7615]),.i2(intermediate_reg_0[7614]),.o(intermediate_reg_1[3807]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7613]),.i2(intermediate_reg_0[7612]),.o(intermediate_reg_1[3806])); 
fsm fsm_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7611]),.i2(intermediate_reg_0[7610]),.o(intermediate_reg_1[3805])); 
fsm fsm_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7609]),.i2(intermediate_reg_0[7608]),.o(intermediate_reg_1[3804])); 
mux_module mux_module_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7607]),.i2(intermediate_reg_0[7606]),.o(intermediate_reg_1[3803]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7605]),.i2(intermediate_reg_0[7604]),.o(intermediate_reg_1[3802]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7603]),.i2(intermediate_reg_0[7602]),.o(intermediate_reg_1[3801])); 
mux_module mux_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7601]),.i2(intermediate_reg_0[7600]),.o(intermediate_reg_1[3800]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7599]),.i2(intermediate_reg_0[7598]),.o(intermediate_reg_1[3799]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7597]),.i2(intermediate_reg_0[7596]),.o(intermediate_reg_1[3798])); 
fsm fsm_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7595]),.i2(intermediate_reg_0[7594]),.o(intermediate_reg_1[3797])); 
mux_module mux_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7593]),.i2(intermediate_reg_0[7592]),.o(intermediate_reg_1[3796]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7591]),.i2(intermediate_reg_0[7590]),.o(intermediate_reg_1[3795])); 
mux_module mux_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7589]),.i2(intermediate_reg_0[7588]),.o(intermediate_reg_1[3794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7587]),.i2(intermediate_reg_0[7586]),.o(intermediate_reg_1[3793]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7585]),.i2(intermediate_reg_0[7584]),.o(intermediate_reg_1[3792]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7583]),.i2(intermediate_reg_0[7582]),.o(intermediate_reg_1[3791]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7581]),.i2(intermediate_reg_0[7580]),.o(intermediate_reg_1[3790])); 
mux_module mux_module_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7579]),.i2(intermediate_reg_0[7578]),.o(intermediate_reg_1[3789]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7577]),.i2(intermediate_reg_0[7576]),.o(intermediate_reg_1[3788]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7575]),.i2(intermediate_reg_0[7574]),.o(intermediate_reg_1[3787]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7573]),.i2(intermediate_reg_0[7572]),.o(intermediate_reg_1[3786]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7571]),.i2(intermediate_reg_0[7570]),.o(intermediate_reg_1[3785]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7569]),.i2(intermediate_reg_0[7568]),.o(intermediate_reg_1[3784]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7567]),.i2(intermediate_reg_0[7566]),.o(intermediate_reg_1[3783])); 
fsm fsm_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7565]),.i2(intermediate_reg_0[7564]),.o(intermediate_reg_1[3782])); 
mux_module mux_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7563]),.i2(intermediate_reg_0[7562]),.o(intermediate_reg_1[3781]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7561]),.i2(intermediate_reg_0[7560]),.o(intermediate_reg_1[3780]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7559]),.i2(intermediate_reg_0[7558]),.o(intermediate_reg_1[3779])); 
fsm fsm_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7557]),.i2(intermediate_reg_0[7556]),.o(intermediate_reg_1[3778])); 
mux_module mux_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7555]),.i2(intermediate_reg_0[7554]),.o(intermediate_reg_1[3777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7553]),.i2(intermediate_reg_0[7552]),.o(intermediate_reg_1[3776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7551]),.i2(intermediate_reg_0[7550]),.o(intermediate_reg_1[3775]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7549]),.i2(intermediate_reg_0[7548]),.o(intermediate_reg_1[3774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7547]),.i2(intermediate_reg_0[7546]),.o(intermediate_reg_1[3773]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7545]),.i2(intermediate_reg_0[7544]),.o(intermediate_reg_1[3772]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7543]),.i2(intermediate_reg_0[7542]),.o(intermediate_reg_1[3771])); 
fsm fsm_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7541]),.i2(intermediate_reg_0[7540]),.o(intermediate_reg_1[3770])); 
mux_module mux_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7539]),.i2(intermediate_reg_0[7538]),.o(intermediate_reg_1[3769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7537]),.i2(intermediate_reg_0[7536]),.o(intermediate_reg_1[3768]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7535]),.i2(intermediate_reg_0[7534]),.o(intermediate_reg_1[3767])); 
mux_module mux_module_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7533]),.i2(intermediate_reg_0[7532]),.o(intermediate_reg_1[3766]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7531]),.i2(intermediate_reg_0[7530]),.o(intermediate_reg_1[3765]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7529]),.i2(intermediate_reg_0[7528]),.o(intermediate_reg_1[3764])); 
mux_module mux_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7527]),.i2(intermediate_reg_0[7526]),.o(intermediate_reg_1[3763]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7525]),.i2(intermediate_reg_0[7524]),.o(intermediate_reg_1[3762]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7523]),.i2(intermediate_reg_0[7522]),.o(intermediate_reg_1[3761]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7521]),.i2(intermediate_reg_0[7520]),.o(intermediate_reg_1[3760])); 
fsm fsm_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7519]),.i2(intermediate_reg_0[7518]),.o(intermediate_reg_1[3759])); 
mux_module mux_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7517]),.i2(intermediate_reg_0[7516]),.o(intermediate_reg_1[3758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7515]),.i2(intermediate_reg_0[7514]),.o(intermediate_reg_1[3757]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7513]),.i2(intermediate_reg_0[7512]),.o(intermediate_reg_1[3756])); 
mux_module mux_module_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7511]),.i2(intermediate_reg_0[7510]),.o(intermediate_reg_1[3755]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7509]),.i2(intermediate_reg_0[7508]),.o(intermediate_reg_1[3754])); 
mux_module mux_module_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7507]),.i2(intermediate_reg_0[7506]),.o(intermediate_reg_1[3753]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7505]),.i2(intermediate_reg_0[7504]),.o(intermediate_reg_1[3752])); 
fsm fsm_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7503]),.i2(intermediate_reg_0[7502]),.o(intermediate_reg_1[3751])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7501]),.i2(intermediate_reg_0[7500]),.o(intermediate_reg_1[3750]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7499]),.i2(intermediate_reg_0[7498]),.o(intermediate_reg_1[3749])); 
fsm fsm_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7497]),.i2(intermediate_reg_0[7496]),.o(intermediate_reg_1[3748])); 
fsm fsm_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7495]),.i2(intermediate_reg_0[7494]),.o(intermediate_reg_1[3747])); 
mux_module mux_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7493]),.i2(intermediate_reg_0[7492]),.o(intermediate_reg_1[3746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7491]),.i2(intermediate_reg_0[7490]),.o(intermediate_reg_1[3745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7489]),.i2(intermediate_reg_0[7488]),.o(intermediate_reg_1[3744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7487]),.i2(intermediate_reg_0[7486]),.o(intermediate_reg_1[3743]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7485]),.i2(intermediate_reg_0[7484]),.o(intermediate_reg_1[3742])); 
fsm fsm_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7483]),.i2(intermediate_reg_0[7482]),.o(intermediate_reg_1[3741])); 
mux_module mux_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7481]),.i2(intermediate_reg_0[7480]),.o(intermediate_reg_1[3740]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7479]),.i2(intermediate_reg_0[7478]),.o(intermediate_reg_1[3739]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7477]),.i2(intermediate_reg_0[7476]),.o(intermediate_reg_1[3738])); 
fsm fsm_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7475]),.i2(intermediate_reg_0[7474]),.o(intermediate_reg_1[3737])); 
mux_module mux_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7473]),.i2(intermediate_reg_0[7472]),.o(intermediate_reg_1[3736]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7471]),.i2(intermediate_reg_0[7470]),.o(intermediate_reg_1[3735])); 
mux_module mux_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7469]),.i2(intermediate_reg_0[7468]),.o(intermediate_reg_1[3734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7467]),.i2(intermediate_reg_0[7466]),.o(intermediate_reg_1[3733]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7465]),.i2(intermediate_reg_0[7464]),.o(intermediate_reg_1[3732]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7463]),.i2(intermediate_reg_0[7462]),.o(intermediate_reg_1[3731])); 
fsm fsm_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7461]),.i2(intermediate_reg_0[7460]),.o(intermediate_reg_1[3730])); 
fsm fsm_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7459]),.i2(intermediate_reg_0[7458]),.o(intermediate_reg_1[3729])); 
mux_module mux_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7457]),.i2(intermediate_reg_0[7456]),.o(intermediate_reg_1[3728]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7455]),.i2(intermediate_reg_0[7454]),.o(intermediate_reg_1[3727]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7453]),.i2(intermediate_reg_0[7452]),.o(intermediate_reg_1[3726]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7451]),.i2(intermediate_reg_0[7450]),.o(intermediate_reg_1[3725])); 
fsm fsm_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7449]),.i2(intermediate_reg_0[7448]),.o(intermediate_reg_1[3724])); 
fsm fsm_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7447]),.i2(intermediate_reg_0[7446]),.o(intermediate_reg_1[3723])); 
fsm fsm_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7445]),.i2(intermediate_reg_0[7444]),.o(intermediate_reg_1[3722])); 
fsm fsm_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7443]),.i2(intermediate_reg_0[7442]),.o(intermediate_reg_1[3721])); 
mux_module mux_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7441]),.i2(intermediate_reg_0[7440]),.o(intermediate_reg_1[3720]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7439]),.i2(intermediate_reg_0[7438]),.o(intermediate_reg_1[3719])); 
fsm fsm_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7437]),.i2(intermediate_reg_0[7436]),.o(intermediate_reg_1[3718])); 
mux_module mux_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7435]),.i2(intermediate_reg_0[7434]),.o(intermediate_reg_1[3717]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7433]),.i2(intermediate_reg_0[7432]),.o(intermediate_reg_1[3716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7431]),.i2(intermediate_reg_0[7430]),.o(intermediate_reg_1[3715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7429]),.i2(intermediate_reg_0[7428]),.o(intermediate_reg_1[3714]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7427]),.i2(intermediate_reg_0[7426]),.o(intermediate_reg_1[3713])); 
fsm fsm_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7425]),.i2(intermediate_reg_0[7424]),.o(intermediate_reg_1[3712])); 
mux_module mux_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7423]),.i2(intermediate_reg_0[7422]),.o(intermediate_reg_1[3711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7421]),.i2(intermediate_reg_0[7420]),.o(intermediate_reg_1[3710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7419]),.i2(intermediate_reg_0[7418]),.o(intermediate_reg_1[3709]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7417]),.i2(intermediate_reg_0[7416]),.o(intermediate_reg_1[3708])); 
fsm fsm_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7415]),.i2(intermediate_reg_0[7414]),.o(intermediate_reg_1[3707])); 
mux_module mux_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7413]),.i2(intermediate_reg_0[7412]),.o(intermediate_reg_1[3706]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7411]),.i2(intermediate_reg_0[7410]),.o(intermediate_reg_1[3705])); 
mux_module mux_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7409]),.i2(intermediate_reg_0[7408]),.o(intermediate_reg_1[3704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7407]),.i2(intermediate_reg_0[7406]),.o(intermediate_reg_1[3703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7405]),.i2(intermediate_reg_0[7404]),.o(intermediate_reg_1[3702]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7403]),.i2(intermediate_reg_0[7402]),.o(intermediate_reg_1[3701]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7401]),.i2(intermediate_reg_0[7400]),.o(intermediate_reg_1[3700]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7399]),.i2(intermediate_reg_0[7398]),.o(intermediate_reg_1[3699]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7397]),.i2(intermediate_reg_0[7396]),.o(intermediate_reg_1[3698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7395]),.i2(intermediate_reg_0[7394]),.o(intermediate_reg_1[3697]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7393]),.i2(intermediate_reg_0[7392]),.o(intermediate_reg_1[3696])); 
mux_module mux_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7391]),.i2(intermediate_reg_0[7390]),.o(intermediate_reg_1[3695]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7389]),.i2(intermediate_reg_0[7388]),.o(intermediate_reg_1[3694])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7387]),.i2(intermediate_reg_0[7386]),.o(intermediate_reg_1[3693]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7385]),.i2(intermediate_reg_0[7384]),.o(intermediate_reg_1[3692])); 
fsm fsm_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7383]),.i2(intermediate_reg_0[7382]),.o(intermediate_reg_1[3691])); 
mux_module mux_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7381]),.i2(intermediate_reg_0[7380]),.o(intermediate_reg_1[3690]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7379]),.i2(intermediate_reg_0[7378]),.o(intermediate_reg_1[3689])); 
fsm fsm_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7377]),.i2(intermediate_reg_0[7376]),.o(intermediate_reg_1[3688])); 
fsm fsm_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7375]),.i2(intermediate_reg_0[7374]),.o(intermediate_reg_1[3687])); 
fsm fsm_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7373]),.i2(intermediate_reg_0[7372]),.o(intermediate_reg_1[3686])); 
fsm fsm_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7371]),.i2(intermediate_reg_0[7370]),.o(intermediate_reg_1[3685])); 
fsm fsm_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7369]),.i2(intermediate_reg_0[7368]),.o(intermediate_reg_1[3684])); 
mux_module mux_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7367]),.i2(intermediate_reg_0[7366]),.o(intermediate_reg_1[3683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7365]),.i2(intermediate_reg_0[7364]),.o(intermediate_reg_1[3682]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7363]),.i2(intermediate_reg_0[7362]),.o(intermediate_reg_1[3681]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7361]),.i2(intermediate_reg_0[7360]),.o(intermediate_reg_1[3680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7359]),.i2(intermediate_reg_0[7358]),.o(intermediate_reg_1[3679]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7357]),.i2(intermediate_reg_0[7356]),.o(intermediate_reg_1[3678])); 
mux_module mux_module_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7355]),.i2(intermediate_reg_0[7354]),.o(intermediate_reg_1[3677]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7353]),.i2(intermediate_reg_0[7352]),.o(intermediate_reg_1[3676])); 
fsm fsm_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7351]),.i2(intermediate_reg_0[7350]),.o(intermediate_reg_1[3675])); 
fsm fsm_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7349]),.i2(intermediate_reg_0[7348]),.o(intermediate_reg_1[3674])); 
fsm fsm_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7347]),.i2(intermediate_reg_0[7346]),.o(intermediate_reg_1[3673])); 
fsm fsm_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7345]),.i2(intermediate_reg_0[7344]),.o(intermediate_reg_1[3672])); 
mux_module mux_module_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7343]),.i2(intermediate_reg_0[7342]),.o(intermediate_reg_1[3671]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7341]),.i2(intermediate_reg_0[7340]),.o(intermediate_reg_1[3670]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7339]),.i2(intermediate_reg_0[7338]),.o(intermediate_reg_1[3669])); 
fsm fsm_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7337]),.i2(intermediate_reg_0[7336]),.o(intermediate_reg_1[3668])); 
fsm fsm_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7335]),.i2(intermediate_reg_0[7334]),.o(intermediate_reg_1[3667])); 
fsm fsm_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7333]),.i2(intermediate_reg_0[7332]),.o(intermediate_reg_1[3666])); 
fsm fsm_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7331]),.i2(intermediate_reg_0[7330]),.o(intermediate_reg_1[3665])); 
fsm fsm_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7329]),.i2(intermediate_reg_0[7328]),.o(intermediate_reg_1[3664])); 
fsm fsm_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7327]),.i2(intermediate_reg_0[7326]),.o(intermediate_reg_1[3663])); 
mux_module mux_module_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7325]),.i2(intermediate_reg_0[7324]),.o(intermediate_reg_1[3662]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7323]),.i2(intermediate_reg_0[7322]),.o(intermediate_reg_1[3661])); 
mux_module mux_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7321]),.i2(intermediate_reg_0[7320]),.o(intermediate_reg_1[3660]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7319]),.i2(intermediate_reg_0[7318]),.o(intermediate_reg_1[3659])); 
mux_module mux_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7317]),.i2(intermediate_reg_0[7316]),.o(intermediate_reg_1[3658]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7315]),.i2(intermediate_reg_0[7314]),.o(intermediate_reg_1[3657])); 
mux_module mux_module_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7313]),.i2(intermediate_reg_0[7312]),.o(intermediate_reg_1[3656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7311]),.i2(intermediate_reg_0[7310]),.o(intermediate_reg_1[3655]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7309]),.i2(intermediate_reg_0[7308]),.o(intermediate_reg_1[3654])); 
mux_module mux_module_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7307]),.i2(intermediate_reg_0[7306]),.o(intermediate_reg_1[3653]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7305]),.i2(intermediate_reg_0[7304]),.o(intermediate_reg_1[3652])); 
fsm fsm_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7303]),.i2(intermediate_reg_0[7302]),.o(intermediate_reg_1[3651])); 
fsm fsm_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7301]),.i2(intermediate_reg_0[7300]),.o(intermediate_reg_1[3650])); 
mux_module mux_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7299]),.i2(intermediate_reg_0[7298]),.o(intermediate_reg_1[3649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7297]),.i2(intermediate_reg_0[7296]),.o(intermediate_reg_1[3648]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7295]),.i2(intermediate_reg_0[7294]),.o(intermediate_reg_1[3647]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7293]),.i2(intermediate_reg_0[7292]),.o(intermediate_reg_1[3646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7291]),.i2(intermediate_reg_0[7290]),.o(intermediate_reg_1[3645]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7289]),.i2(intermediate_reg_0[7288]),.o(intermediate_reg_1[3644]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7287]),.i2(intermediate_reg_0[7286]),.o(intermediate_reg_1[3643]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7285]),.i2(intermediate_reg_0[7284]),.o(intermediate_reg_1[3642])); 
mux_module mux_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7283]),.i2(intermediate_reg_0[7282]),.o(intermediate_reg_1[3641]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7281]),.i2(intermediate_reg_0[7280]),.o(intermediate_reg_1[3640])); 
mux_module mux_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7279]),.i2(intermediate_reg_0[7278]),.o(intermediate_reg_1[3639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7277]),.i2(intermediate_reg_0[7276]),.o(intermediate_reg_1[3638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7275]),.i2(intermediate_reg_0[7274]),.o(intermediate_reg_1[3637])); 
fsm fsm_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7273]),.i2(intermediate_reg_0[7272]),.o(intermediate_reg_1[3636])); 
mux_module mux_module_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7271]),.i2(intermediate_reg_0[7270]),.o(intermediate_reg_1[3635]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7269]),.i2(intermediate_reg_0[7268]),.o(intermediate_reg_1[3634])); 
fsm fsm_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7267]),.i2(intermediate_reg_0[7266]),.o(intermediate_reg_1[3633])); 
mux_module mux_module_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7265]),.i2(intermediate_reg_0[7264]),.o(intermediate_reg_1[3632]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7263]),.i2(intermediate_reg_0[7262]),.o(intermediate_reg_1[3631])); 
fsm fsm_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7261]),.i2(intermediate_reg_0[7260]),.o(intermediate_reg_1[3630])); 
fsm fsm_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7259]),.i2(intermediate_reg_0[7258]),.o(intermediate_reg_1[3629])); 
fsm fsm_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7257]),.i2(intermediate_reg_0[7256]),.o(intermediate_reg_1[3628])); 
mux_module mux_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7255]),.i2(intermediate_reg_0[7254]),.o(intermediate_reg_1[3627]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7253]),.i2(intermediate_reg_0[7252]),.o(intermediate_reg_1[3626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7251]),.i2(intermediate_reg_0[7250]),.o(intermediate_reg_1[3625])); 
mux_module mux_module_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7249]),.i2(intermediate_reg_0[7248]),.o(intermediate_reg_1[3624]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7247]),.i2(intermediate_reg_0[7246]),.o(intermediate_reg_1[3623]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7245]),.i2(intermediate_reg_0[7244]),.o(intermediate_reg_1[3622]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7243]),.i2(intermediate_reg_0[7242]),.o(intermediate_reg_1[3621])); 
mux_module mux_module_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7241]),.i2(intermediate_reg_0[7240]),.o(intermediate_reg_1[3620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7239]),.i2(intermediate_reg_0[7238]),.o(intermediate_reg_1[3619]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7237]),.i2(intermediate_reg_0[7236]),.o(intermediate_reg_1[3618]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7235]),.i2(intermediate_reg_0[7234]),.o(intermediate_reg_1[3617]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7233]),.i2(intermediate_reg_0[7232]),.o(intermediate_reg_1[3616])); 
mux_module mux_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7231]),.i2(intermediate_reg_0[7230]),.o(intermediate_reg_1[3615]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7229]),.i2(intermediate_reg_0[7228]),.o(intermediate_reg_1[3614])); 
mux_module mux_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7227]),.i2(intermediate_reg_0[7226]),.o(intermediate_reg_1[3613]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7225]),.i2(intermediate_reg_0[7224]),.o(intermediate_reg_1[3612])); 
fsm fsm_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7223]),.i2(intermediate_reg_0[7222]),.o(intermediate_reg_1[3611])); 
mux_module mux_module_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7221]),.i2(intermediate_reg_0[7220]),.o(intermediate_reg_1[3610]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7219]),.i2(intermediate_reg_0[7218]),.o(intermediate_reg_1[3609])); 
mux_module mux_module_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7217]),.i2(intermediate_reg_0[7216]),.o(intermediate_reg_1[3608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7215]),.i2(intermediate_reg_0[7214]),.o(intermediate_reg_1[3607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7213]),.i2(intermediate_reg_0[7212]),.o(intermediate_reg_1[3606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7211]),.i2(intermediate_reg_0[7210]),.o(intermediate_reg_1[3605]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7209]),.i2(intermediate_reg_0[7208]),.o(intermediate_reg_1[3604])); 
fsm fsm_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7207]),.i2(intermediate_reg_0[7206]),.o(intermediate_reg_1[3603])); 
fsm fsm_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7205]),.i2(intermediate_reg_0[7204]),.o(intermediate_reg_1[3602])); 
mux_module mux_module_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7203]),.i2(intermediate_reg_0[7202]),.o(intermediate_reg_1[3601]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7201]),.i2(intermediate_reg_0[7200]),.o(intermediate_reg_1[3600])); 
mux_module mux_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7199]),.i2(intermediate_reg_0[7198]),.o(intermediate_reg_1[3599]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7197]),.i2(intermediate_reg_0[7196]),.o(intermediate_reg_1[3598])); 
fsm fsm_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7195]),.i2(intermediate_reg_0[7194]),.o(intermediate_reg_1[3597])); 
mux_module mux_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7193]),.i2(intermediate_reg_0[7192]),.o(intermediate_reg_1[3596]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7191]),.i2(intermediate_reg_0[7190]),.o(intermediate_reg_1[3595]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7189]),.i2(intermediate_reg_0[7188]),.o(intermediate_reg_1[3594])); 
fsm fsm_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7187]),.i2(intermediate_reg_0[7186]),.o(intermediate_reg_1[3593])); 
fsm fsm_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7185]),.i2(intermediate_reg_0[7184]),.o(intermediate_reg_1[3592])); 
fsm fsm_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7183]),.i2(intermediate_reg_0[7182]),.o(intermediate_reg_1[3591])); 
mux_module mux_module_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7181]),.i2(intermediate_reg_0[7180]),.o(intermediate_reg_1[3590]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7179]),.i2(intermediate_reg_0[7178]),.o(intermediate_reg_1[3589]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7177]),.i2(intermediate_reg_0[7176]),.o(intermediate_reg_1[3588]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7175]),.i2(intermediate_reg_0[7174]),.o(intermediate_reg_1[3587])); 
fsm fsm_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7173]),.i2(intermediate_reg_0[7172]),.o(intermediate_reg_1[3586])); 
fsm fsm_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7171]),.i2(intermediate_reg_0[7170]),.o(intermediate_reg_1[3585])); 
mux_module mux_module_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7169]),.i2(intermediate_reg_0[7168]),.o(intermediate_reg_1[3584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7167]),.i2(intermediate_reg_0[7166]),.o(intermediate_reg_1[3583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7165]),.i2(intermediate_reg_0[7164]),.o(intermediate_reg_1[3582]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7163]),.i2(intermediate_reg_0[7162]),.o(intermediate_reg_1[3581]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7161]),.i2(intermediate_reg_0[7160]),.o(intermediate_reg_1[3580])); 
fsm fsm_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7159]),.i2(intermediate_reg_0[7158]),.o(intermediate_reg_1[3579])); 
mux_module mux_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7157]),.i2(intermediate_reg_0[7156]),.o(intermediate_reg_1[3578]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7155]),.i2(intermediate_reg_0[7154]),.o(intermediate_reg_1[3577])); 
fsm fsm_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7153]),.i2(intermediate_reg_0[7152]),.o(intermediate_reg_1[3576])); 
mux_module mux_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7151]),.i2(intermediate_reg_0[7150]),.o(intermediate_reg_1[3575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7149]),.i2(intermediate_reg_0[7148]),.o(intermediate_reg_1[3574]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7147]),.i2(intermediate_reg_0[7146]),.o(intermediate_reg_1[3573]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7145]),.i2(intermediate_reg_0[7144]),.o(intermediate_reg_1[3572])); 
fsm fsm_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7143]),.i2(intermediate_reg_0[7142]),.o(intermediate_reg_1[3571])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7141]),.i2(intermediate_reg_0[7140]),.o(intermediate_reg_1[3570]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7139]),.i2(intermediate_reg_0[7138]),.o(intermediate_reg_1[3569])); 
fsm fsm_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7137]),.i2(intermediate_reg_0[7136]),.o(intermediate_reg_1[3568])); 
fsm fsm_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7135]),.i2(intermediate_reg_0[7134]),.o(intermediate_reg_1[3567])); 
fsm fsm_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7133]),.i2(intermediate_reg_0[7132]),.o(intermediate_reg_1[3566])); 
mux_module mux_module_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7131]),.i2(intermediate_reg_0[7130]),.o(intermediate_reg_1[3565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7129]),.i2(intermediate_reg_0[7128]),.o(intermediate_reg_1[3564]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7127]),.i2(intermediate_reg_0[7126]),.o(intermediate_reg_1[3563])); 
mux_module mux_module_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7125]),.i2(intermediate_reg_0[7124]),.o(intermediate_reg_1[3562]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7123]),.i2(intermediate_reg_0[7122]),.o(intermediate_reg_1[3561])); 
fsm fsm_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7121]),.i2(intermediate_reg_0[7120]),.o(intermediate_reg_1[3560])); 
fsm fsm_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7119]),.i2(intermediate_reg_0[7118]),.o(intermediate_reg_1[3559])); 
fsm fsm_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7117]),.i2(intermediate_reg_0[7116]),.o(intermediate_reg_1[3558])); 
fsm fsm_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7115]),.i2(intermediate_reg_0[7114]),.o(intermediate_reg_1[3557])); 
mux_module mux_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7113]),.i2(intermediate_reg_0[7112]),.o(intermediate_reg_1[3556]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7111]),.i2(intermediate_reg_0[7110]),.o(intermediate_reg_1[3555])); 
mux_module mux_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7109]),.i2(intermediate_reg_0[7108]),.o(intermediate_reg_1[3554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7107]),.i2(intermediate_reg_0[7106]),.o(intermediate_reg_1[3553]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7105]),.i2(intermediate_reg_0[7104]),.o(intermediate_reg_1[3552])); 
fsm fsm_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7103]),.i2(intermediate_reg_0[7102]),.o(intermediate_reg_1[3551])); 
mux_module mux_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7101]),.i2(intermediate_reg_0[7100]),.o(intermediate_reg_1[3550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7099]),.i2(intermediate_reg_0[7098]),.o(intermediate_reg_1[3549]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7097]),.i2(intermediate_reg_0[7096]),.o(intermediate_reg_1[3548])); 
mux_module mux_module_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7095]),.i2(intermediate_reg_0[7094]),.o(intermediate_reg_1[3547]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7093]),.i2(intermediate_reg_0[7092]),.o(intermediate_reg_1[3546])); 
mux_module mux_module_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7091]),.i2(intermediate_reg_0[7090]),.o(intermediate_reg_1[3545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7089]),.i2(intermediate_reg_0[7088]),.o(intermediate_reg_1[3544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7087]),.i2(intermediate_reg_0[7086]),.o(intermediate_reg_1[3543]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7085]),.i2(intermediate_reg_0[7084]),.o(intermediate_reg_1[3542])); 
mux_module mux_module_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7083]),.i2(intermediate_reg_0[7082]),.o(intermediate_reg_1[3541]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7081]),.i2(intermediate_reg_0[7080]),.o(intermediate_reg_1[3540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7079]),.i2(intermediate_reg_0[7078]),.o(intermediate_reg_1[3539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7077]),.i2(intermediate_reg_0[7076]),.o(intermediate_reg_1[3538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7075]),.i2(intermediate_reg_0[7074]),.o(intermediate_reg_1[3537]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7073]),.i2(intermediate_reg_0[7072]),.o(intermediate_reg_1[3536]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7071]),.i2(intermediate_reg_0[7070]),.o(intermediate_reg_1[3535]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7069]),.i2(intermediate_reg_0[7068]),.o(intermediate_reg_1[3534]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7067]),.i2(intermediate_reg_0[7066]),.o(intermediate_reg_1[3533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7065]),.i2(intermediate_reg_0[7064]),.o(intermediate_reg_1[3532]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7063]),.i2(intermediate_reg_0[7062]),.o(intermediate_reg_1[3531])); 
fsm fsm_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7061]),.i2(intermediate_reg_0[7060]),.o(intermediate_reg_1[3530])); 
fsm fsm_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7059]),.i2(intermediate_reg_0[7058]),.o(intermediate_reg_1[3529])); 
fsm fsm_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7057]),.i2(intermediate_reg_0[7056]),.o(intermediate_reg_1[3528])); 
mux_module mux_module_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7055]),.i2(intermediate_reg_0[7054]),.o(intermediate_reg_1[3527]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7053]),.i2(intermediate_reg_0[7052]),.o(intermediate_reg_1[3526])); 
mux_module mux_module_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7051]),.i2(intermediate_reg_0[7050]),.o(intermediate_reg_1[3525]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7049]),.i2(intermediate_reg_0[7048]),.o(intermediate_reg_1[3524])); 
fsm fsm_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7047]),.i2(intermediate_reg_0[7046]),.o(intermediate_reg_1[3523])); 
fsm fsm_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7045]),.i2(intermediate_reg_0[7044]),.o(intermediate_reg_1[3522])); 
fsm fsm_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7043]),.i2(intermediate_reg_0[7042]),.o(intermediate_reg_1[3521])); 
fsm fsm_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7041]),.i2(intermediate_reg_0[7040]),.o(intermediate_reg_1[3520])); 
mux_module mux_module_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7039]),.i2(intermediate_reg_0[7038]),.o(intermediate_reg_1[3519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7037]),.i2(intermediate_reg_0[7036]),.o(intermediate_reg_1[3518]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7035]),.i2(intermediate_reg_0[7034]),.o(intermediate_reg_1[3517]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7033]),.i2(intermediate_reg_0[7032]),.o(intermediate_reg_1[3516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7031]),.i2(intermediate_reg_0[7030]),.o(intermediate_reg_1[3515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7029]),.i2(intermediate_reg_0[7028]),.o(intermediate_reg_1[3514]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7027]),.i2(intermediate_reg_0[7026]),.o(intermediate_reg_1[3513]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7025]),.i2(intermediate_reg_0[7024]),.o(intermediate_reg_1[3512])); 
fsm fsm_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7023]),.i2(intermediate_reg_0[7022]),.o(intermediate_reg_1[3511])); 
fsm fsm_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7021]),.i2(intermediate_reg_0[7020]),.o(intermediate_reg_1[3510])); 
mux_module mux_module_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7019]),.i2(intermediate_reg_0[7018]),.o(intermediate_reg_1[3509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7017]),.i2(intermediate_reg_0[7016]),.o(intermediate_reg_1[3508]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7015]),.i2(intermediate_reg_0[7014]),.o(intermediate_reg_1[3507])); 
mux_module mux_module_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7013]),.i2(intermediate_reg_0[7012]),.o(intermediate_reg_1[3506]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7011]),.i2(intermediate_reg_0[7010]),.o(intermediate_reg_1[3505])); 
mux_module mux_module_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7009]),.i2(intermediate_reg_0[7008]),.o(intermediate_reg_1[3504]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7007]),.i2(intermediate_reg_0[7006]),.o(intermediate_reg_1[3503]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7005]),.i2(intermediate_reg_0[7004]),.o(intermediate_reg_1[3502])); 
fsm fsm_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7003]),.i2(intermediate_reg_0[7002]),.o(intermediate_reg_1[3501])); 
fsm fsm_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7001]),.i2(intermediate_reg_0[7000]),.o(intermediate_reg_1[3500])); 
fsm fsm_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6999]),.i2(intermediate_reg_0[6998]),.o(intermediate_reg_1[3499])); 
fsm fsm_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6997]),.i2(intermediate_reg_0[6996]),.o(intermediate_reg_1[3498])); 
mux_module mux_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6995]),.i2(intermediate_reg_0[6994]),.o(intermediate_reg_1[3497]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6993]),.i2(intermediate_reg_0[6992]),.o(intermediate_reg_1[3496])); 
mux_module mux_module_inst_1_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6991]),.i2(intermediate_reg_0[6990]),.o(intermediate_reg_1[3495]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6989]),.i2(intermediate_reg_0[6988]),.o(intermediate_reg_1[3494]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6987]),.i2(intermediate_reg_0[6986]),.o(intermediate_reg_1[3493])); 
fsm fsm_inst_1_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6985]),.i2(intermediate_reg_0[6984]),.o(intermediate_reg_1[3492])); 
fsm fsm_inst_1_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6983]),.i2(intermediate_reg_0[6982]),.o(intermediate_reg_1[3491])); 
mux_module mux_module_inst_1_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6981]),.i2(intermediate_reg_0[6980]),.o(intermediate_reg_1[3490]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6979]),.i2(intermediate_reg_0[6978]),.o(intermediate_reg_1[3489]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6977]),.i2(intermediate_reg_0[6976]),.o(intermediate_reg_1[3488])); 
fsm fsm_inst_1_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6975]),.i2(intermediate_reg_0[6974]),.o(intermediate_reg_1[3487])); 
fsm fsm_inst_1_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6973]),.i2(intermediate_reg_0[6972]),.o(intermediate_reg_1[3486])); 
fsm fsm_inst_1_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6971]),.i2(intermediate_reg_0[6970]),.o(intermediate_reg_1[3485])); 
mux_module mux_module_inst_1_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6969]),.i2(intermediate_reg_0[6968]),.o(intermediate_reg_1[3484]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6967]),.i2(intermediate_reg_0[6966]),.o(intermediate_reg_1[3483])); 
fsm fsm_inst_1_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6965]),.i2(intermediate_reg_0[6964]),.o(intermediate_reg_1[3482])); 
fsm fsm_inst_1_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6963]),.i2(intermediate_reg_0[6962]),.o(intermediate_reg_1[3481])); 
fsm fsm_inst_1_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6961]),.i2(intermediate_reg_0[6960]),.o(intermediate_reg_1[3480])); 
mux_module mux_module_inst_1_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6959]),.i2(intermediate_reg_0[6958]),.o(intermediate_reg_1[3479]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6957]),.i2(intermediate_reg_0[6956]),.o(intermediate_reg_1[3478]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6955]),.i2(intermediate_reg_0[6954]),.o(intermediate_reg_1[3477]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6953]),.i2(intermediate_reg_0[6952]),.o(intermediate_reg_1[3476])); 
mux_module mux_module_inst_1_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6951]),.i2(intermediate_reg_0[6950]),.o(intermediate_reg_1[3475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6949]),.i2(intermediate_reg_0[6948]),.o(intermediate_reg_1[3474]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6947]),.i2(intermediate_reg_0[6946]),.o(intermediate_reg_1[3473])); 
fsm fsm_inst_1_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6945]),.i2(intermediate_reg_0[6944]),.o(intermediate_reg_1[3472])); 
fsm fsm_inst_1_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6943]),.i2(intermediate_reg_0[6942]),.o(intermediate_reg_1[3471])); 
mux_module mux_module_inst_1_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6941]),.i2(intermediate_reg_0[6940]),.o(intermediate_reg_1[3470]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6939]),.i2(intermediate_reg_0[6938]),.o(intermediate_reg_1[3469]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6937]),.i2(intermediate_reg_0[6936]),.o(intermediate_reg_1[3468]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6935]),.i2(intermediate_reg_0[6934]),.o(intermediate_reg_1[3467])); 
mux_module mux_module_inst_1_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6933]),.i2(intermediate_reg_0[6932]),.o(intermediate_reg_1[3466]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6931]),.i2(intermediate_reg_0[6930]),.o(intermediate_reg_1[3465])); 
mux_module mux_module_inst_1_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6929]),.i2(intermediate_reg_0[6928]),.o(intermediate_reg_1[3464]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6927]),.i2(intermediate_reg_0[6926]),.o(intermediate_reg_1[3463])); 
fsm fsm_inst_1_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6925]),.i2(intermediate_reg_0[6924]),.o(intermediate_reg_1[3462])); 
fsm fsm_inst_1_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6923]),.i2(intermediate_reg_0[6922]),.o(intermediate_reg_1[3461])); 
fsm fsm_inst_1_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6921]),.i2(intermediate_reg_0[6920]),.o(intermediate_reg_1[3460])); 
mux_module mux_module_inst_1_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6919]),.i2(intermediate_reg_0[6918]),.o(intermediate_reg_1[3459]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6917]),.i2(intermediate_reg_0[6916]),.o(intermediate_reg_1[3458])); 
fsm fsm_inst_1_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6915]),.i2(intermediate_reg_0[6914]),.o(intermediate_reg_1[3457])); 
mux_module mux_module_inst_1_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6913]),.i2(intermediate_reg_0[6912]),.o(intermediate_reg_1[3456]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6911]),.i2(intermediate_reg_0[6910]),.o(intermediate_reg_1[3455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6909]),.i2(intermediate_reg_0[6908]),.o(intermediate_reg_1[3454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6907]),.i2(intermediate_reg_0[6906]),.o(intermediate_reg_1[3453]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6905]),.i2(intermediate_reg_0[6904]),.o(intermediate_reg_1[3452])); 
mux_module mux_module_inst_1_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6903]),.i2(intermediate_reg_0[6902]),.o(intermediate_reg_1[3451]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6901]),.i2(intermediate_reg_0[6900]),.o(intermediate_reg_1[3450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6899]),.i2(intermediate_reg_0[6898]),.o(intermediate_reg_1[3449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6897]),.i2(intermediate_reg_0[6896]),.o(intermediate_reg_1[3448])); 
mux_module mux_module_inst_1_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6895]),.i2(intermediate_reg_0[6894]),.o(intermediate_reg_1[3447]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6893]),.i2(intermediate_reg_0[6892]),.o(intermediate_reg_1[3446]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6891]),.i2(intermediate_reg_0[6890]),.o(intermediate_reg_1[3445]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6889]),.i2(intermediate_reg_0[6888]),.o(intermediate_reg_1[3444]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6887]),.i2(intermediate_reg_0[6886]),.o(intermediate_reg_1[3443])); 
mux_module mux_module_inst_1_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6885]),.i2(intermediate_reg_0[6884]),.o(intermediate_reg_1[3442]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6883]),.i2(intermediate_reg_0[6882]),.o(intermediate_reg_1[3441])); 
fsm fsm_inst_1_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6881]),.i2(intermediate_reg_0[6880]),.o(intermediate_reg_1[3440])); 
mux_module mux_module_inst_1_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6879]),.i2(intermediate_reg_0[6878]),.o(intermediate_reg_1[3439]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6877]),.i2(intermediate_reg_0[6876]),.o(intermediate_reg_1[3438])); 
mux_module mux_module_inst_1_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6875]),.i2(intermediate_reg_0[6874]),.o(intermediate_reg_1[3437]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6873]),.i2(intermediate_reg_0[6872]),.o(intermediate_reg_1[3436]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6871]),.i2(intermediate_reg_0[6870]),.o(intermediate_reg_1[3435])); 
mux_module mux_module_inst_1_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6869]),.i2(intermediate_reg_0[6868]),.o(intermediate_reg_1[3434]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6867]),.i2(intermediate_reg_0[6866]),.o(intermediate_reg_1[3433])); 
fsm fsm_inst_1_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6865]),.i2(intermediate_reg_0[6864]),.o(intermediate_reg_1[3432])); 
fsm fsm_inst_1_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6863]),.i2(intermediate_reg_0[6862]),.o(intermediate_reg_1[3431])); 
mux_module mux_module_inst_1_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6861]),.i2(intermediate_reg_0[6860]),.o(intermediate_reg_1[3430]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6859]),.i2(intermediate_reg_0[6858]),.o(intermediate_reg_1[3429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6857]),.i2(intermediate_reg_0[6856]),.o(intermediate_reg_1[3428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6855]),.i2(intermediate_reg_0[6854]),.o(intermediate_reg_1[3427]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6853]),.i2(intermediate_reg_0[6852]),.o(intermediate_reg_1[3426]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6851]),.i2(intermediate_reg_0[6850]),.o(intermediate_reg_1[3425])); 
fsm fsm_inst_1_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6849]),.i2(intermediate_reg_0[6848]),.o(intermediate_reg_1[3424])); 
fsm fsm_inst_1_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6847]),.i2(intermediate_reg_0[6846]),.o(intermediate_reg_1[3423])); 
mux_module mux_module_inst_1_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6845]),.i2(intermediate_reg_0[6844]),.o(intermediate_reg_1[3422]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6843]),.i2(intermediate_reg_0[6842]),.o(intermediate_reg_1[3421])); 
fsm fsm_inst_1_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6841]),.i2(intermediate_reg_0[6840]),.o(intermediate_reg_1[3420])); 
fsm fsm_inst_1_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6839]),.i2(intermediate_reg_0[6838]),.o(intermediate_reg_1[3419])); 
mux_module mux_module_inst_1_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6837]),.i2(intermediate_reg_0[6836]),.o(intermediate_reg_1[3418]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6835]),.i2(intermediate_reg_0[6834]),.o(intermediate_reg_1[3417])); 
mux_module mux_module_inst_1_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6833]),.i2(intermediate_reg_0[6832]),.o(intermediate_reg_1[3416]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6831]),.i2(intermediate_reg_0[6830]),.o(intermediate_reg_1[3415])); 
mux_module mux_module_inst_1_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6829]),.i2(intermediate_reg_0[6828]),.o(intermediate_reg_1[3414]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6827]),.i2(intermediate_reg_0[6826]),.o(intermediate_reg_1[3413])); 
mux_module mux_module_inst_1_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6825]),.i2(intermediate_reg_0[6824]),.o(intermediate_reg_1[3412]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6823]),.i2(intermediate_reg_0[6822]),.o(intermediate_reg_1[3411])); 
mux_module mux_module_inst_1_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6821]),.i2(intermediate_reg_0[6820]),.o(intermediate_reg_1[3410]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6819]),.i2(intermediate_reg_0[6818]),.o(intermediate_reg_1[3409])); 
fsm fsm_inst_1_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6817]),.i2(intermediate_reg_0[6816]),.o(intermediate_reg_1[3408])); 
fsm fsm_inst_1_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6815]),.i2(intermediate_reg_0[6814]),.o(intermediate_reg_1[3407])); 
fsm fsm_inst_1_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6813]),.i2(intermediate_reg_0[6812]),.o(intermediate_reg_1[3406])); 
fsm fsm_inst_1_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6811]),.i2(intermediate_reg_0[6810]),.o(intermediate_reg_1[3405])); 
mux_module mux_module_inst_1_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6809]),.i2(intermediate_reg_0[6808]),.o(intermediate_reg_1[3404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6807]),.i2(intermediate_reg_0[6806]),.o(intermediate_reg_1[3403])); 
mux_module mux_module_inst_1_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6805]),.i2(intermediate_reg_0[6804]),.o(intermediate_reg_1[3402]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6803]),.i2(intermediate_reg_0[6802]),.o(intermediate_reg_1[3401]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6801]),.i2(intermediate_reg_0[6800]),.o(intermediate_reg_1[3400])); 
fsm fsm_inst_1_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6799]),.i2(intermediate_reg_0[6798]),.o(intermediate_reg_1[3399])); 
mux_module mux_module_inst_1_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6797]),.i2(intermediate_reg_0[6796]),.o(intermediate_reg_1[3398]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6795]),.i2(intermediate_reg_0[6794]),.o(intermediate_reg_1[3397]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6793]),.i2(intermediate_reg_0[6792]),.o(intermediate_reg_1[3396])); 
fsm fsm_inst_1_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6791]),.i2(intermediate_reg_0[6790]),.o(intermediate_reg_1[3395])); 
mux_module mux_module_inst_1_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6789]),.i2(intermediate_reg_0[6788]),.o(intermediate_reg_1[3394]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6787]),.i2(intermediate_reg_0[6786]),.o(intermediate_reg_1[3393])); 
fsm fsm_inst_1_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6785]),.i2(intermediate_reg_0[6784]),.o(intermediate_reg_1[3392])); 
mux_module mux_module_inst_1_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6783]),.i2(intermediate_reg_0[6782]),.o(intermediate_reg_1[3391]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6781]),.i2(intermediate_reg_0[6780]),.o(intermediate_reg_1[3390]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6779]),.i2(intermediate_reg_0[6778]),.o(intermediate_reg_1[3389]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6777]),.i2(intermediate_reg_0[6776]),.o(intermediate_reg_1[3388]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6775]),.i2(intermediate_reg_0[6774]),.o(intermediate_reg_1[3387])); 
fsm fsm_inst_1_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6773]),.i2(intermediate_reg_0[6772]),.o(intermediate_reg_1[3386])); 
fsm fsm_inst_1_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6771]),.i2(intermediate_reg_0[6770]),.o(intermediate_reg_1[3385])); 
mux_module mux_module_inst_1_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6769]),.i2(intermediate_reg_0[6768]),.o(intermediate_reg_1[3384]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6767]),.i2(intermediate_reg_0[6766]),.o(intermediate_reg_1[3383])); 
fsm fsm_inst_1_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6765]),.i2(intermediate_reg_0[6764]),.o(intermediate_reg_1[3382])); 
fsm fsm_inst_1_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6763]),.i2(intermediate_reg_0[6762]),.o(intermediate_reg_1[3381])); 
mux_module mux_module_inst_1_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6761]),.i2(intermediate_reg_0[6760]),.o(intermediate_reg_1[3380]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6759]),.i2(intermediate_reg_0[6758]),.o(intermediate_reg_1[3379])); 
mux_module mux_module_inst_1_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6757]),.i2(intermediate_reg_0[6756]),.o(intermediate_reg_1[3378]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6755]),.i2(intermediate_reg_0[6754]),.o(intermediate_reg_1[3377])); 
mux_module mux_module_inst_1_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6753]),.i2(intermediate_reg_0[6752]),.o(intermediate_reg_1[3376]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6751]),.i2(intermediate_reg_0[6750]),.o(intermediate_reg_1[3375])); 
mux_module mux_module_inst_1_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6749]),.i2(intermediate_reg_0[6748]),.o(intermediate_reg_1[3374]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6747]),.i2(intermediate_reg_0[6746]),.o(intermediate_reg_1[3373])); 
mux_module mux_module_inst_1_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6745]),.i2(intermediate_reg_0[6744]),.o(intermediate_reg_1[3372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6743]),.i2(intermediate_reg_0[6742]),.o(intermediate_reg_1[3371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6741]),.i2(intermediate_reg_0[6740]),.o(intermediate_reg_1[3370]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6739]),.i2(intermediate_reg_0[6738]),.o(intermediate_reg_1[3369]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6737]),.i2(intermediate_reg_0[6736]),.o(intermediate_reg_1[3368])); 
fsm fsm_inst_1_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6735]),.i2(intermediate_reg_0[6734]),.o(intermediate_reg_1[3367])); 
mux_module mux_module_inst_1_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6733]),.i2(intermediate_reg_0[6732]),.o(intermediate_reg_1[3366]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6731]),.i2(intermediate_reg_0[6730]),.o(intermediate_reg_1[3365])); 
fsm fsm_inst_1_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6729]),.i2(intermediate_reg_0[6728]),.o(intermediate_reg_1[3364])); 
fsm fsm_inst_1_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6727]),.i2(intermediate_reg_0[6726]),.o(intermediate_reg_1[3363])); 
fsm fsm_inst_1_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6725]),.i2(intermediate_reg_0[6724]),.o(intermediate_reg_1[3362])); 
fsm fsm_inst_1_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6723]),.i2(intermediate_reg_0[6722]),.o(intermediate_reg_1[3361])); 
fsm fsm_inst_1_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6721]),.i2(intermediate_reg_0[6720]),.o(intermediate_reg_1[3360])); 
fsm fsm_inst_1_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6719]),.i2(intermediate_reg_0[6718]),.o(intermediate_reg_1[3359])); 
fsm fsm_inst_1_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6717]),.i2(intermediate_reg_0[6716]),.o(intermediate_reg_1[3358])); 
fsm fsm_inst_1_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6715]),.i2(intermediate_reg_0[6714]),.o(intermediate_reg_1[3357])); 
mux_module mux_module_inst_1_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6713]),.i2(intermediate_reg_0[6712]),.o(intermediate_reg_1[3356]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6711]),.i2(intermediate_reg_0[6710]),.o(intermediate_reg_1[3355])); 
mux_module mux_module_inst_1_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6709]),.i2(intermediate_reg_0[6708]),.o(intermediate_reg_1[3354]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6707]),.i2(intermediate_reg_0[6706]),.o(intermediate_reg_1[3353])); 
fsm fsm_inst_1_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6705]),.i2(intermediate_reg_0[6704]),.o(intermediate_reg_1[3352])); 
fsm fsm_inst_1_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6703]),.i2(intermediate_reg_0[6702]),.o(intermediate_reg_1[3351])); 
fsm fsm_inst_1_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6701]),.i2(intermediate_reg_0[6700]),.o(intermediate_reg_1[3350])); 
fsm fsm_inst_1_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6699]),.i2(intermediate_reg_0[6698]),.o(intermediate_reg_1[3349])); 
mux_module mux_module_inst_1_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6697]),.i2(intermediate_reg_0[6696]),.o(intermediate_reg_1[3348]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6695]),.i2(intermediate_reg_0[6694]),.o(intermediate_reg_1[3347]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6693]),.i2(intermediate_reg_0[6692]),.o(intermediate_reg_1[3346])); 
mux_module mux_module_inst_1_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6691]),.i2(intermediate_reg_0[6690]),.o(intermediate_reg_1[3345]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6689]),.i2(intermediate_reg_0[6688]),.o(intermediate_reg_1[3344])); 
fsm fsm_inst_1_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6687]),.i2(intermediate_reg_0[6686]),.o(intermediate_reg_1[3343])); 
mux_module mux_module_inst_1_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6685]),.i2(intermediate_reg_0[6684]),.o(intermediate_reg_1[3342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6683]),.i2(intermediate_reg_0[6682]),.o(intermediate_reg_1[3341]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6681]),.i2(intermediate_reg_0[6680]),.o(intermediate_reg_1[3340])); 
mux_module mux_module_inst_1_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6679]),.i2(intermediate_reg_0[6678]),.o(intermediate_reg_1[3339]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6677]),.i2(intermediate_reg_0[6676]),.o(intermediate_reg_1[3338]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6675]),.i2(intermediate_reg_0[6674]),.o(intermediate_reg_1[3337])); 
mux_module mux_module_inst_1_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6673]),.i2(intermediate_reg_0[6672]),.o(intermediate_reg_1[3336]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6671]),.i2(intermediate_reg_0[6670]),.o(intermediate_reg_1[3335]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6669]),.i2(intermediate_reg_0[6668]),.o(intermediate_reg_1[3334]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6667]),.i2(intermediate_reg_0[6666]),.o(intermediate_reg_1[3333])); 
fsm fsm_inst_1_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6665]),.i2(intermediate_reg_0[6664]),.o(intermediate_reg_1[3332])); 
mux_module mux_module_inst_1_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6663]),.i2(intermediate_reg_0[6662]),.o(intermediate_reg_1[3331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6661]),.i2(intermediate_reg_0[6660]),.o(intermediate_reg_1[3330]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6659]),.i2(intermediate_reg_0[6658]),.o(intermediate_reg_1[3329])); 
fsm fsm_inst_1_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6657]),.i2(intermediate_reg_0[6656]),.o(intermediate_reg_1[3328])); 
fsm fsm_inst_1_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6655]),.i2(intermediate_reg_0[6654]),.o(intermediate_reg_1[3327])); 
mux_module mux_module_inst_1_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6653]),.i2(intermediate_reg_0[6652]),.o(intermediate_reg_1[3326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6651]),.i2(intermediate_reg_0[6650]),.o(intermediate_reg_1[3325]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6649]),.i2(intermediate_reg_0[6648]),.o(intermediate_reg_1[3324])); 
mux_module mux_module_inst_1_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6647]),.i2(intermediate_reg_0[6646]),.o(intermediate_reg_1[3323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6645]),.i2(intermediate_reg_0[6644]),.o(intermediate_reg_1[3322]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6643]),.i2(intermediate_reg_0[6642]),.o(intermediate_reg_1[3321])); 
mux_module mux_module_inst_1_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6641]),.i2(intermediate_reg_0[6640]),.o(intermediate_reg_1[3320]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6639]),.i2(intermediate_reg_0[6638]),.o(intermediate_reg_1[3319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6637]),.i2(intermediate_reg_0[6636]),.o(intermediate_reg_1[3318]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6635]),.i2(intermediate_reg_0[6634]),.o(intermediate_reg_1[3317])); 
fsm fsm_inst_1_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6633]),.i2(intermediate_reg_0[6632]),.o(intermediate_reg_1[3316])); 
fsm fsm_inst_1_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6631]),.i2(intermediate_reg_0[6630]),.o(intermediate_reg_1[3315])); 
fsm fsm_inst_1_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6629]),.i2(intermediate_reg_0[6628]),.o(intermediate_reg_1[3314])); 
mux_module mux_module_inst_1_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6627]),.i2(intermediate_reg_0[6626]),.o(intermediate_reg_1[3313]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6625]),.i2(intermediate_reg_0[6624]),.o(intermediate_reg_1[3312])); 
mux_module mux_module_inst_1_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6623]),.i2(intermediate_reg_0[6622]),.o(intermediate_reg_1[3311]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6621]),.i2(intermediate_reg_0[6620]),.o(intermediate_reg_1[3310])); 
mux_module mux_module_inst_1_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6619]),.i2(intermediate_reg_0[6618]),.o(intermediate_reg_1[3309]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6617]),.i2(intermediate_reg_0[6616]),.o(intermediate_reg_1[3308])); 
fsm fsm_inst_1_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6615]),.i2(intermediate_reg_0[6614]),.o(intermediate_reg_1[3307])); 
fsm fsm_inst_1_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6613]),.i2(intermediate_reg_0[6612]),.o(intermediate_reg_1[3306])); 
fsm fsm_inst_1_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6611]),.i2(intermediate_reg_0[6610]),.o(intermediate_reg_1[3305])); 
fsm fsm_inst_1_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6609]),.i2(intermediate_reg_0[6608]),.o(intermediate_reg_1[3304])); 
mux_module mux_module_inst_1_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6607]),.i2(intermediate_reg_0[6606]),.o(intermediate_reg_1[3303]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6605]),.i2(intermediate_reg_0[6604]),.o(intermediate_reg_1[3302])); 
fsm fsm_inst_1_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6603]),.i2(intermediate_reg_0[6602]),.o(intermediate_reg_1[3301])); 
mux_module mux_module_inst_1_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6601]),.i2(intermediate_reg_0[6600]),.o(intermediate_reg_1[3300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6599]),.i2(intermediate_reg_0[6598]),.o(intermediate_reg_1[3299]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6597]),.i2(intermediate_reg_0[6596]),.o(intermediate_reg_1[3298])); 
mux_module mux_module_inst_1_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6595]),.i2(intermediate_reg_0[6594]),.o(intermediate_reg_1[3297]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6593]),.i2(intermediate_reg_0[6592]),.o(intermediate_reg_1[3296])); 
fsm fsm_inst_1_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6591]),.i2(intermediate_reg_0[6590]),.o(intermediate_reg_1[3295])); 
fsm fsm_inst_1_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6589]),.i2(intermediate_reg_0[6588]),.o(intermediate_reg_1[3294])); 
mux_module mux_module_inst_1_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6587]),.i2(intermediate_reg_0[6586]),.o(intermediate_reg_1[3293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6585]),.i2(intermediate_reg_0[6584]),.o(intermediate_reg_1[3292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6583]),.i2(intermediate_reg_0[6582]),.o(intermediate_reg_1[3291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6581]),.i2(intermediate_reg_0[6580]),.o(intermediate_reg_1[3290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6579]),.i2(intermediate_reg_0[6578]),.o(intermediate_reg_1[3289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6577]),.i2(intermediate_reg_0[6576]),.o(intermediate_reg_1[3288]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6575]),.i2(intermediate_reg_0[6574]),.o(intermediate_reg_1[3287])); 
fsm fsm_inst_1_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6573]),.i2(intermediate_reg_0[6572]),.o(intermediate_reg_1[3286])); 
fsm fsm_inst_1_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6571]),.i2(intermediate_reg_0[6570]),.o(intermediate_reg_1[3285])); 
fsm fsm_inst_1_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6569]),.i2(intermediate_reg_0[6568]),.o(intermediate_reg_1[3284])); 
fsm fsm_inst_1_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6567]),.i2(intermediate_reg_0[6566]),.o(intermediate_reg_1[3283])); 
fsm fsm_inst_1_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6565]),.i2(intermediate_reg_0[6564]),.o(intermediate_reg_1[3282])); 
mux_module mux_module_inst_1_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6563]),.i2(intermediate_reg_0[6562]),.o(intermediate_reg_1[3281]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6561]),.i2(intermediate_reg_0[6560]),.o(intermediate_reg_1[3280])); 
fsm fsm_inst_1_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6559]),.i2(intermediate_reg_0[6558]),.o(intermediate_reg_1[3279])); 
mux_module mux_module_inst_1_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6557]),.i2(intermediate_reg_0[6556]),.o(intermediate_reg_1[3278]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6555]),.i2(intermediate_reg_0[6554]),.o(intermediate_reg_1[3277])); 
fsm fsm_inst_1_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6553]),.i2(intermediate_reg_0[6552]),.o(intermediate_reg_1[3276])); 
mux_module mux_module_inst_1_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6551]),.i2(intermediate_reg_0[6550]),.o(intermediate_reg_1[3275]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6549]),.i2(intermediate_reg_0[6548]),.o(intermediate_reg_1[3274])); 
mux_module mux_module_inst_1_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6547]),.i2(intermediate_reg_0[6546]),.o(intermediate_reg_1[3273]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6545]),.i2(intermediate_reg_0[6544]),.o(intermediate_reg_1[3272])); 
mux_module mux_module_inst_1_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6543]),.i2(intermediate_reg_0[6542]),.o(intermediate_reg_1[3271]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6541]),.i2(intermediate_reg_0[6540]),.o(intermediate_reg_1[3270]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6539]),.i2(intermediate_reg_0[6538]),.o(intermediate_reg_1[3269])); 
fsm fsm_inst_1_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6537]),.i2(intermediate_reg_0[6536]),.o(intermediate_reg_1[3268])); 
mux_module mux_module_inst_1_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6535]),.i2(intermediate_reg_0[6534]),.o(intermediate_reg_1[3267]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6533]),.i2(intermediate_reg_0[6532]),.o(intermediate_reg_1[3266])); 
fsm fsm_inst_1_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6531]),.i2(intermediate_reg_0[6530]),.o(intermediate_reg_1[3265])); 
fsm fsm_inst_1_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6529]),.i2(intermediate_reg_0[6528]),.o(intermediate_reg_1[3264])); 
fsm fsm_inst_1_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6527]),.i2(intermediate_reg_0[6526]),.o(intermediate_reg_1[3263])); 
fsm fsm_inst_1_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6525]),.i2(intermediate_reg_0[6524]),.o(intermediate_reg_1[3262])); 
mux_module mux_module_inst_1_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6523]),.i2(intermediate_reg_0[6522]),.o(intermediate_reg_1[3261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6521]),.i2(intermediate_reg_0[6520]),.o(intermediate_reg_1[3260]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6519]),.i2(intermediate_reg_0[6518]),.o(intermediate_reg_1[3259])); 
fsm fsm_inst_1_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6517]),.i2(intermediate_reg_0[6516]),.o(intermediate_reg_1[3258])); 
fsm fsm_inst_1_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6515]),.i2(intermediate_reg_0[6514]),.o(intermediate_reg_1[3257])); 
mux_module mux_module_inst_1_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6513]),.i2(intermediate_reg_0[6512]),.o(intermediate_reg_1[3256]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6511]),.i2(intermediate_reg_0[6510]),.o(intermediate_reg_1[3255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6509]),.i2(intermediate_reg_0[6508]),.o(intermediate_reg_1[3254]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6507]),.i2(intermediate_reg_0[6506]),.o(intermediate_reg_1[3253])); 
mux_module mux_module_inst_1_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6505]),.i2(intermediate_reg_0[6504]),.o(intermediate_reg_1[3252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6503]),.i2(intermediate_reg_0[6502]),.o(intermediate_reg_1[3251]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6501]),.i2(intermediate_reg_0[6500]),.o(intermediate_reg_1[3250])); 
mux_module mux_module_inst_1_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6499]),.i2(intermediate_reg_0[6498]),.o(intermediate_reg_1[3249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6497]),.i2(intermediate_reg_0[6496]),.o(intermediate_reg_1[3248]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6495]),.i2(intermediate_reg_0[6494]),.o(intermediate_reg_1[3247])); 
fsm fsm_inst_1_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6493]),.i2(intermediate_reg_0[6492]),.o(intermediate_reg_1[3246])); 
fsm fsm_inst_1_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6491]),.i2(intermediate_reg_0[6490]),.o(intermediate_reg_1[3245])); 
fsm fsm_inst_1_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6489]),.i2(intermediate_reg_0[6488]),.o(intermediate_reg_1[3244])); 
fsm fsm_inst_1_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6487]),.i2(intermediate_reg_0[6486]),.o(intermediate_reg_1[3243])); 
mux_module mux_module_inst_1_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6485]),.i2(intermediate_reg_0[6484]),.o(intermediate_reg_1[3242]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6483]),.i2(intermediate_reg_0[6482]),.o(intermediate_reg_1[3241]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6481]),.i2(intermediate_reg_0[6480]),.o(intermediate_reg_1[3240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6479]),.i2(intermediate_reg_0[6478]),.o(intermediate_reg_1[3239]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6477]),.i2(intermediate_reg_0[6476]),.o(intermediate_reg_1[3238])); 
mux_module mux_module_inst_1_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6475]),.i2(intermediate_reg_0[6474]),.o(intermediate_reg_1[3237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6473]),.i2(intermediate_reg_0[6472]),.o(intermediate_reg_1[3236]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6471]),.i2(intermediate_reg_0[6470]),.o(intermediate_reg_1[3235])); 
fsm fsm_inst_1_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6469]),.i2(intermediate_reg_0[6468]),.o(intermediate_reg_1[3234])); 
mux_module mux_module_inst_1_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6467]),.i2(intermediate_reg_0[6466]),.o(intermediate_reg_1[3233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6465]),.i2(intermediate_reg_0[6464]),.o(intermediate_reg_1[3232]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6463]),.i2(intermediate_reg_0[6462]),.o(intermediate_reg_1[3231])); 
fsm fsm_inst_1_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6461]),.i2(intermediate_reg_0[6460]),.o(intermediate_reg_1[3230])); 
fsm fsm_inst_1_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6459]),.i2(intermediate_reg_0[6458]),.o(intermediate_reg_1[3229])); 
fsm fsm_inst_1_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6457]),.i2(intermediate_reg_0[6456]),.o(intermediate_reg_1[3228])); 
mux_module mux_module_inst_1_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6455]),.i2(intermediate_reg_0[6454]),.o(intermediate_reg_1[3227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6453]),.i2(intermediate_reg_0[6452]),.o(intermediate_reg_1[3226]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6451]),.i2(intermediate_reg_0[6450]),.o(intermediate_reg_1[3225]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6449]),.i2(intermediate_reg_0[6448]),.o(intermediate_reg_1[3224])); 
fsm fsm_inst_1_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6447]),.i2(intermediate_reg_0[6446]),.o(intermediate_reg_1[3223])); 
fsm fsm_inst_1_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6445]),.i2(intermediate_reg_0[6444]),.o(intermediate_reg_1[3222])); 
fsm fsm_inst_1_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6443]),.i2(intermediate_reg_0[6442]),.o(intermediate_reg_1[3221])); 
mux_module mux_module_inst_1_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6441]),.i2(intermediate_reg_0[6440]),.o(intermediate_reg_1[3220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6439]),.i2(intermediate_reg_0[6438]),.o(intermediate_reg_1[3219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6437]),.i2(intermediate_reg_0[6436]),.o(intermediate_reg_1[3218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6435]),.i2(intermediate_reg_0[6434]),.o(intermediate_reg_1[3217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6433]),.i2(intermediate_reg_0[6432]),.o(intermediate_reg_1[3216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6431]),.i2(intermediate_reg_0[6430]),.o(intermediate_reg_1[3215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6429]),.i2(intermediate_reg_0[6428]),.o(intermediate_reg_1[3214]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6427]),.i2(intermediate_reg_0[6426]),.o(intermediate_reg_1[3213])); 
mux_module mux_module_inst_1_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6425]),.i2(intermediate_reg_0[6424]),.o(intermediate_reg_1[3212]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6423]),.i2(intermediate_reg_0[6422]),.o(intermediate_reg_1[3211])); 
mux_module mux_module_inst_1_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6421]),.i2(intermediate_reg_0[6420]),.o(intermediate_reg_1[3210]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6419]),.i2(intermediate_reg_0[6418]),.o(intermediate_reg_1[3209]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6417]),.i2(intermediate_reg_0[6416]),.o(intermediate_reg_1[3208])); 
mux_module mux_module_inst_1_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6415]),.i2(intermediate_reg_0[6414]),.o(intermediate_reg_1[3207]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6413]),.i2(intermediate_reg_0[6412]),.o(intermediate_reg_1[3206])); 
fsm fsm_inst_1_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6411]),.i2(intermediate_reg_0[6410]),.o(intermediate_reg_1[3205])); 
fsm fsm_inst_1_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6409]),.i2(intermediate_reg_0[6408]),.o(intermediate_reg_1[3204])); 
fsm fsm_inst_1_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6407]),.i2(intermediate_reg_0[6406]),.o(intermediate_reg_1[3203])); 
mux_module mux_module_inst_1_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6405]),.i2(intermediate_reg_0[6404]),.o(intermediate_reg_1[3202]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6403]),.i2(intermediate_reg_0[6402]),.o(intermediate_reg_1[3201])); 
mux_module mux_module_inst_1_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6401]),.i2(intermediate_reg_0[6400]),.o(intermediate_reg_1[3200]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6399]),.i2(intermediate_reg_0[6398]),.o(intermediate_reg_1[3199])); 
fsm fsm_inst_1_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6397]),.i2(intermediate_reg_0[6396]),.o(intermediate_reg_1[3198])); 
fsm fsm_inst_1_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6395]),.i2(intermediate_reg_0[6394]),.o(intermediate_reg_1[3197])); 
mux_module mux_module_inst_1_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6393]),.i2(intermediate_reg_0[6392]),.o(intermediate_reg_1[3196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6391]),.i2(intermediate_reg_0[6390]),.o(intermediate_reg_1[3195]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6389]),.i2(intermediate_reg_0[6388]),.o(intermediate_reg_1[3194])); 
mux_module mux_module_inst_1_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6387]),.i2(intermediate_reg_0[6386]),.o(intermediate_reg_1[3193]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6385]),.i2(intermediate_reg_0[6384]),.o(intermediate_reg_1[3192])); 
fsm fsm_inst_1_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6383]),.i2(intermediate_reg_0[6382]),.o(intermediate_reg_1[3191])); 
fsm fsm_inst_1_1649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6381]),.i2(intermediate_reg_0[6380]),.o(intermediate_reg_1[3190])); 
fsm fsm_inst_1_1650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6379]),.i2(intermediate_reg_0[6378]),.o(intermediate_reg_1[3189])); 
mux_module mux_module_inst_1_1651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6377]),.i2(intermediate_reg_0[6376]),.o(intermediate_reg_1[3188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6375]),.i2(intermediate_reg_0[6374]),.o(intermediate_reg_1[3187]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6373]),.i2(intermediate_reg_0[6372]),.o(intermediate_reg_1[3186])); 
fsm fsm_inst_1_1654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6371]),.i2(intermediate_reg_0[6370]),.o(intermediate_reg_1[3185])); 
mux_module mux_module_inst_1_1655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6369]),.i2(intermediate_reg_0[6368]),.o(intermediate_reg_1[3184]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6367]),.i2(intermediate_reg_0[6366]),.o(intermediate_reg_1[3183])); 
mux_module mux_module_inst_1_1657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6365]),.i2(intermediate_reg_0[6364]),.o(intermediate_reg_1[3182]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6363]),.i2(intermediate_reg_0[6362]),.o(intermediate_reg_1[3181])); 
mux_module mux_module_inst_1_1659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6361]),.i2(intermediate_reg_0[6360]),.o(intermediate_reg_1[3180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6359]),.i2(intermediate_reg_0[6358]),.o(intermediate_reg_1[3179]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6357]),.i2(intermediate_reg_0[6356]),.o(intermediate_reg_1[3178])); 
fsm fsm_inst_1_1662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6355]),.i2(intermediate_reg_0[6354]),.o(intermediate_reg_1[3177])); 
fsm fsm_inst_1_1663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6353]),.i2(intermediate_reg_0[6352]),.o(intermediate_reg_1[3176])); 
mux_module mux_module_inst_1_1664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6351]),.i2(intermediate_reg_0[6350]),.o(intermediate_reg_1[3175]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6349]),.i2(intermediate_reg_0[6348]),.o(intermediate_reg_1[3174])); 
mux_module mux_module_inst_1_1666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6347]),.i2(intermediate_reg_0[6346]),.o(intermediate_reg_1[3173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6345]),.i2(intermediate_reg_0[6344]),.o(intermediate_reg_1[3172]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6343]),.i2(intermediate_reg_0[6342]),.o(intermediate_reg_1[3171])); 
fsm fsm_inst_1_1669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6341]),.i2(intermediate_reg_0[6340]),.o(intermediate_reg_1[3170])); 
mux_module mux_module_inst_1_1670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6339]),.i2(intermediate_reg_0[6338]),.o(intermediate_reg_1[3169]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6337]),.i2(intermediate_reg_0[6336]),.o(intermediate_reg_1[3168])); 
mux_module mux_module_inst_1_1672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6335]),.i2(intermediate_reg_0[6334]),.o(intermediate_reg_1[3167]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6333]),.i2(intermediate_reg_0[6332]),.o(intermediate_reg_1[3166]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6331]),.i2(intermediate_reg_0[6330]),.o(intermediate_reg_1[3165])); 
mux_module mux_module_inst_1_1675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6329]),.i2(intermediate_reg_0[6328]),.o(intermediate_reg_1[3164]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6327]),.i2(intermediate_reg_0[6326]),.o(intermediate_reg_1[3163])); 
mux_module mux_module_inst_1_1677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6325]),.i2(intermediate_reg_0[6324]),.o(intermediate_reg_1[3162]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6323]),.i2(intermediate_reg_0[6322]),.o(intermediate_reg_1[3161])); 
mux_module mux_module_inst_1_1679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6321]),.i2(intermediate_reg_0[6320]),.o(intermediate_reg_1[3160]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6319]),.i2(intermediate_reg_0[6318]),.o(intermediate_reg_1[3159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6317]),.i2(intermediate_reg_0[6316]),.o(intermediate_reg_1[3158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6315]),.i2(intermediate_reg_0[6314]),.o(intermediate_reg_1[3157]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6313]),.i2(intermediate_reg_0[6312]),.o(intermediate_reg_1[3156]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6311]),.i2(intermediate_reg_0[6310]),.o(intermediate_reg_1[3155]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6309]),.i2(intermediate_reg_0[6308]),.o(intermediate_reg_1[3154])); 
mux_module mux_module_inst_1_1686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6307]),.i2(intermediate_reg_0[6306]),.o(intermediate_reg_1[3153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6305]),.i2(intermediate_reg_0[6304]),.o(intermediate_reg_1[3152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6303]),.i2(intermediate_reg_0[6302]),.o(intermediate_reg_1[3151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6301]),.i2(intermediate_reg_0[6300]),.o(intermediate_reg_1[3150]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6299]),.i2(intermediate_reg_0[6298]),.o(intermediate_reg_1[3149])); 
fsm fsm_inst_1_1691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6297]),.i2(intermediate_reg_0[6296]),.o(intermediate_reg_1[3148])); 
mux_module mux_module_inst_1_1692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6295]),.i2(intermediate_reg_0[6294]),.o(intermediate_reg_1[3147]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6293]),.i2(intermediate_reg_0[6292]),.o(intermediate_reg_1[3146])); 
mux_module mux_module_inst_1_1694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6291]),.i2(intermediate_reg_0[6290]),.o(intermediate_reg_1[3145]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6289]),.i2(intermediate_reg_0[6288]),.o(intermediate_reg_1[3144])); 
fsm fsm_inst_1_1696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6287]),.i2(intermediate_reg_0[6286]),.o(intermediate_reg_1[3143])); 
mux_module mux_module_inst_1_1697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6285]),.i2(intermediate_reg_0[6284]),.o(intermediate_reg_1[3142]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6283]),.i2(intermediate_reg_0[6282]),.o(intermediate_reg_1[3141]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6281]),.i2(intermediate_reg_0[6280]),.o(intermediate_reg_1[3140])); 
fsm fsm_inst_1_1700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6279]),.i2(intermediate_reg_0[6278]),.o(intermediate_reg_1[3139])); 
fsm fsm_inst_1_1701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6277]),.i2(intermediate_reg_0[6276]),.o(intermediate_reg_1[3138])); 
fsm fsm_inst_1_1702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6275]),.i2(intermediate_reg_0[6274]),.o(intermediate_reg_1[3137])); 
fsm fsm_inst_1_1703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6273]),.i2(intermediate_reg_0[6272]),.o(intermediate_reg_1[3136])); 
mux_module mux_module_inst_1_1704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6271]),.i2(intermediate_reg_0[6270]),.o(intermediate_reg_1[3135]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6269]),.i2(intermediate_reg_0[6268]),.o(intermediate_reg_1[3134]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6267]),.i2(intermediate_reg_0[6266]),.o(intermediate_reg_1[3133])); 
fsm fsm_inst_1_1707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6265]),.i2(intermediate_reg_0[6264]),.o(intermediate_reg_1[3132])); 
fsm fsm_inst_1_1708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6263]),.i2(intermediate_reg_0[6262]),.o(intermediate_reg_1[3131])); 
fsm fsm_inst_1_1709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6261]),.i2(intermediate_reg_0[6260]),.o(intermediate_reg_1[3130])); 
fsm fsm_inst_1_1710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6259]),.i2(intermediate_reg_0[6258]),.o(intermediate_reg_1[3129])); 
fsm fsm_inst_1_1711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6257]),.i2(intermediate_reg_0[6256]),.o(intermediate_reg_1[3128])); 
mux_module mux_module_inst_1_1712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6255]),.i2(intermediate_reg_0[6254]),.o(intermediate_reg_1[3127]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6253]),.i2(intermediate_reg_0[6252]),.o(intermediate_reg_1[3126])); 
fsm fsm_inst_1_1714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6251]),.i2(intermediate_reg_0[6250]),.o(intermediate_reg_1[3125])); 
fsm fsm_inst_1_1715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6249]),.i2(intermediate_reg_0[6248]),.o(intermediate_reg_1[3124])); 
fsm fsm_inst_1_1716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6247]),.i2(intermediate_reg_0[6246]),.o(intermediate_reg_1[3123])); 
mux_module mux_module_inst_1_1717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6245]),.i2(intermediate_reg_0[6244]),.o(intermediate_reg_1[3122]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6243]),.i2(intermediate_reg_0[6242]),.o(intermediate_reg_1[3121])); 
fsm fsm_inst_1_1719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6241]),.i2(intermediate_reg_0[6240]),.o(intermediate_reg_1[3120])); 
fsm fsm_inst_1_1720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6239]),.i2(intermediate_reg_0[6238]),.o(intermediate_reg_1[3119])); 
fsm fsm_inst_1_1721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6237]),.i2(intermediate_reg_0[6236]),.o(intermediate_reg_1[3118])); 
fsm fsm_inst_1_1722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6235]),.i2(intermediate_reg_0[6234]),.o(intermediate_reg_1[3117])); 
mux_module mux_module_inst_1_1723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6233]),.i2(intermediate_reg_0[6232]),.o(intermediate_reg_1[3116]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6231]),.i2(intermediate_reg_0[6230]),.o(intermediate_reg_1[3115])); 
fsm fsm_inst_1_1725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6229]),.i2(intermediate_reg_0[6228]),.o(intermediate_reg_1[3114])); 
fsm fsm_inst_1_1726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6227]),.i2(intermediate_reg_0[6226]),.o(intermediate_reg_1[3113])); 
mux_module mux_module_inst_1_1727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6225]),.i2(intermediate_reg_0[6224]),.o(intermediate_reg_1[3112]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6223]),.i2(intermediate_reg_0[6222]),.o(intermediate_reg_1[3111])); 
fsm fsm_inst_1_1729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6221]),.i2(intermediate_reg_0[6220]),.o(intermediate_reg_1[3110])); 
mux_module mux_module_inst_1_1730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6219]),.i2(intermediate_reg_0[6218]),.o(intermediate_reg_1[3109]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6217]),.i2(intermediate_reg_0[6216]),.o(intermediate_reg_1[3108])); 
fsm fsm_inst_1_1732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6215]),.i2(intermediate_reg_0[6214]),.o(intermediate_reg_1[3107])); 
fsm fsm_inst_1_1733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6213]),.i2(intermediate_reg_0[6212]),.o(intermediate_reg_1[3106])); 
fsm fsm_inst_1_1734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6211]),.i2(intermediate_reg_0[6210]),.o(intermediate_reg_1[3105])); 
mux_module mux_module_inst_1_1735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6209]),.i2(intermediate_reg_0[6208]),.o(intermediate_reg_1[3104]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6207]),.i2(intermediate_reg_0[6206]),.o(intermediate_reg_1[3103])); 
fsm fsm_inst_1_1737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6205]),.i2(intermediate_reg_0[6204]),.o(intermediate_reg_1[3102])); 
fsm fsm_inst_1_1738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6203]),.i2(intermediate_reg_0[6202]),.o(intermediate_reg_1[3101])); 
mux_module mux_module_inst_1_1739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6201]),.i2(intermediate_reg_0[6200]),.o(intermediate_reg_1[3100]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6199]),.i2(intermediate_reg_0[6198]),.o(intermediate_reg_1[3099])); 
mux_module mux_module_inst_1_1741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6197]),.i2(intermediate_reg_0[6196]),.o(intermediate_reg_1[3098]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6195]),.i2(intermediate_reg_0[6194]),.o(intermediate_reg_1[3097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6193]),.i2(intermediate_reg_0[6192]),.o(intermediate_reg_1[3096]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6191]),.i2(intermediate_reg_0[6190]),.o(intermediate_reg_1[3095])); 
mux_module mux_module_inst_1_1745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6189]),.i2(intermediate_reg_0[6188]),.o(intermediate_reg_1[3094]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6187]),.i2(intermediate_reg_0[6186]),.o(intermediate_reg_1[3093])); 
mux_module mux_module_inst_1_1747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6185]),.i2(intermediate_reg_0[6184]),.o(intermediate_reg_1[3092]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6183]),.i2(intermediate_reg_0[6182]),.o(intermediate_reg_1[3091]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6181]),.i2(intermediate_reg_0[6180]),.o(intermediate_reg_1[3090])); 
fsm fsm_inst_1_1750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6179]),.i2(intermediate_reg_0[6178]),.o(intermediate_reg_1[3089])); 
fsm fsm_inst_1_1751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6177]),.i2(intermediate_reg_0[6176]),.o(intermediate_reg_1[3088])); 
mux_module mux_module_inst_1_1752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6175]),.i2(intermediate_reg_0[6174]),.o(intermediate_reg_1[3087]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6173]),.i2(intermediate_reg_0[6172]),.o(intermediate_reg_1[3086])); 
mux_module mux_module_inst_1_1754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6171]),.i2(intermediate_reg_0[6170]),.o(intermediate_reg_1[3085]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6169]),.i2(intermediate_reg_0[6168]),.o(intermediate_reg_1[3084]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6167]),.i2(intermediate_reg_0[6166]),.o(intermediate_reg_1[3083])); 
mux_module mux_module_inst_1_1757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6165]),.i2(intermediate_reg_0[6164]),.o(intermediate_reg_1[3082]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6163]),.i2(intermediate_reg_0[6162]),.o(intermediate_reg_1[3081]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6161]),.i2(intermediate_reg_0[6160]),.o(intermediate_reg_1[3080])); 
mux_module mux_module_inst_1_1760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6159]),.i2(intermediate_reg_0[6158]),.o(intermediate_reg_1[3079]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6157]),.i2(intermediate_reg_0[6156]),.o(intermediate_reg_1[3078]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6155]),.i2(intermediate_reg_0[6154]),.o(intermediate_reg_1[3077]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6153]),.i2(intermediate_reg_0[6152]),.o(intermediate_reg_1[3076]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6151]),.i2(intermediate_reg_0[6150]),.o(intermediate_reg_1[3075])); 
fsm fsm_inst_1_1765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6149]),.i2(intermediate_reg_0[6148]),.o(intermediate_reg_1[3074])); 
mux_module mux_module_inst_1_1766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6147]),.i2(intermediate_reg_0[6146]),.o(intermediate_reg_1[3073]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6145]),.i2(intermediate_reg_0[6144]),.o(intermediate_reg_1[3072])); 
mux_module mux_module_inst_1_1768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6143]),.i2(intermediate_reg_0[6142]),.o(intermediate_reg_1[3071]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6141]),.i2(intermediate_reg_0[6140]),.o(intermediate_reg_1[3070]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6139]),.i2(intermediate_reg_0[6138]),.o(intermediate_reg_1[3069])); 
mux_module mux_module_inst_1_1771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6137]),.i2(intermediate_reg_0[6136]),.o(intermediate_reg_1[3068]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6135]),.i2(intermediate_reg_0[6134]),.o(intermediate_reg_1[3067])); 
fsm fsm_inst_1_1773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6133]),.i2(intermediate_reg_0[6132]),.o(intermediate_reg_1[3066])); 
mux_module mux_module_inst_1_1774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6131]),.i2(intermediate_reg_0[6130]),.o(intermediate_reg_1[3065]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6129]),.i2(intermediate_reg_0[6128]),.o(intermediate_reg_1[3064]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6127]),.i2(intermediate_reg_0[6126]),.o(intermediate_reg_1[3063])); 
fsm fsm_inst_1_1777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6125]),.i2(intermediate_reg_0[6124]),.o(intermediate_reg_1[3062])); 
fsm fsm_inst_1_1778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6123]),.i2(intermediate_reg_0[6122]),.o(intermediate_reg_1[3061])); 
mux_module mux_module_inst_1_1779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6121]),.i2(intermediate_reg_0[6120]),.o(intermediate_reg_1[3060]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6119]),.i2(intermediate_reg_0[6118]),.o(intermediate_reg_1[3059]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6117]),.i2(intermediate_reg_0[6116]),.o(intermediate_reg_1[3058])); 
mux_module mux_module_inst_1_1782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6115]),.i2(intermediate_reg_0[6114]),.o(intermediate_reg_1[3057]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6113]),.i2(intermediate_reg_0[6112]),.o(intermediate_reg_1[3056])); 
mux_module mux_module_inst_1_1784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6111]),.i2(intermediate_reg_0[6110]),.o(intermediate_reg_1[3055]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6109]),.i2(intermediate_reg_0[6108]),.o(intermediate_reg_1[3054]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6107]),.i2(intermediate_reg_0[6106]),.o(intermediate_reg_1[3053]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6105]),.i2(intermediate_reg_0[6104]),.o(intermediate_reg_1[3052]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6103]),.i2(intermediate_reg_0[6102]),.o(intermediate_reg_1[3051]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6101]),.i2(intermediate_reg_0[6100]),.o(intermediate_reg_1[3050])); 
mux_module mux_module_inst_1_1790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6099]),.i2(intermediate_reg_0[6098]),.o(intermediate_reg_1[3049]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6097]),.i2(intermediate_reg_0[6096]),.o(intermediate_reg_1[3048])); 
fsm fsm_inst_1_1792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6095]),.i2(intermediate_reg_0[6094]),.o(intermediate_reg_1[3047])); 
mux_module mux_module_inst_1_1793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6093]),.i2(intermediate_reg_0[6092]),.o(intermediate_reg_1[3046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6091]),.i2(intermediate_reg_0[6090]),.o(intermediate_reg_1[3045]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6089]),.i2(intermediate_reg_0[6088]),.o(intermediate_reg_1[3044]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6087]),.i2(intermediate_reg_0[6086]),.o(intermediate_reg_1[3043])); 
mux_module mux_module_inst_1_1797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6085]),.i2(intermediate_reg_0[6084]),.o(intermediate_reg_1[3042]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6083]),.i2(intermediate_reg_0[6082]),.o(intermediate_reg_1[3041])); 
fsm fsm_inst_1_1799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6081]),.i2(intermediate_reg_0[6080]),.o(intermediate_reg_1[3040])); 
mux_module mux_module_inst_1_1800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6079]),.i2(intermediate_reg_0[6078]),.o(intermediate_reg_1[3039]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6077]),.i2(intermediate_reg_0[6076]),.o(intermediate_reg_1[3038]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6075]),.i2(intermediate_reg_0[6074]),.o(intermediate_reg_1[3037]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6073]),.i2(intermediate_reg_0[6072]),.o(intermediate_reg_1[3036])); 
mux_module mux_module_inst_1_1804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6071]),.i2(intermediate_reg_0[6070]),.o(intermediate_reg_1[3035]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6069]),.i2(intermediate_reg_0[6068]),.o(intermediate_reg_1[3034]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6067]),.i2(intermediate_reg_0[6066]),.o(intermediate_reg_1[3033]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6065]),.i2(intermediate_reg_0[6064]),.o(intermediate_reg_1[3032])); 
fsm fsm_inst_1_1808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6063]),.i2(intermediate_reg_0[6062]),.o(intermediate_reg_1[3031])); 
fsm fsm_inst_1_1809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6061]),.i2(intermediate_reg_0[6060]),.o(intermediate_reg_1[3030])); 
mux_module mux_module_inst_1_1810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6059]),.i2(intermediate_reg_0[6058]),.o(intermediate_reg_1[3029]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6057]),.i2(intermediate_reg_0[6056]),.o(intermediate_reg_1[3028])); 
fsm fsm_inst_1_1812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6055]),.i2(intermediate_reg_0[6054]),.o(intermediate_reg_1[3027])); 
fsm fsm_inst_1_1813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6053]),.i2(intermediate_reg_0[6052]),.o(intermediate_reg_1[3026])); 
mux_module mux_module_inst_1_1814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6051]),.i2(intermediate_reg_0[6050]),.o(intermediate_reg_1[3025]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6049]),.i2(intermediate_reg_0[6048]),.o(intermediate_reg_1[3024])); 
fsm fsm_inst_1_1816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6047]),.i2(intermediate_reg_0[6046]),.o(intermediate_reg_1[3023])); 
mux_module mux_module_inst_1_1817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6045]),.i2(intermediate_reg_0[6044]),.o(intermediate_reg_1[3022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6043]),.i2(intermediate_reg_0[6042]),.o(intermediate_reg_1[3021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6041]),.i2(intermediate_reg_0[6040]),.o(intermediate_reg_1[3020]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6039]),.i2(intermediate_reg_0[6038]),.o(intermediate_reg_1[3019])); 
fsm fsm_inst_1_1821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6037]),.i2(intermediate_reg_0[6036]),.o(intermediate_reg_1[3018])); 
mux_module mux_module_inst_1_1822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6035]),.i2(intermediate_reg_0[6034]),.o(intermediate_reg_1[3017]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6033]),.i2(intermediate_reg_0[6032]),.o(intermediate_reg_1[3016]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6031]),.i2(intermediate_reg_0[6030]),.o(intermediate_reg_1[3015])); 
mux_module mux_module_inst_1_1825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6029]),.i2(intermediate_reg_0[6028]),.o(intermediate_reg_1[3014]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6027]),.i2(intermediate_reg_0[6026]),.o(intermediate_reg_1[3013]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6025]),.i2(intermediate_reg_0[6024]),.o(intermediate_reg_1[3012]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6023]),.i2(intermediate_reg_0[6022]),.o(intermediate_reg_1[3011]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6021]),.i2(intermediate_reg_0[6020]),.o(intermediate_reg_1[3010]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6019]),.i2(intermediate_reg_0[6018]),.o(intermediate_reg_1[3009]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6017]),.i2(intermediate_reg_0[6016]),.o(intermediate_reg_1[3008]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6015]),.i2(intermediate_reg_0[6014]),.o(intermediate_reg_1[3007]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6013]),.i2(intermediate_reg_0[6012]),.o(intermediate_reg_1[3006]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6011]),.i2(intermediate_reg_0[6010]),.o(intermediate_reg_1[3005])); 
mux_module mux_module_inst_1_1835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6009]),.i2(intermediate_reg_0[6008]),.o(intermediate_reg_1[3004]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6007]),.i2(intermediate_reg_0[6006]),.o(intermediate_reg_1[3003]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6005]),.i2(intermediate_reg_0[6004]),.o(intermediate_reg_1[3002]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6003]),.i2(intermediate_reg_0[6002]),.o(intermediate_reg_1[3001])); 
mux_module mux_module_inst_1_1839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[6001]),.i2(intermediate_reg_0[6000]),.o(intermediate_reg_1[3000]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5999]),.i2(intermediate_reg_0[5998]),.o(intermediate_reg_1[2999]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5997]),.i2(intermediate_reg_0[5996]),.o(intermediate_reg_1[2998]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5995]),.i2(intermediate_reg_0[5994]),.o(intermediate_reg_1[2997])); 
fsm fsm_inst_1_1843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5993]),.i2(intermediate_reg_0[5992]),.o(intermediate_reg_1[2996])); 
fsm fsm_inst_1_1844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5991]),.i2(intermediate_reg_0[5990]),.o(intermediate_reg_1[2995])); 
mux_module mux_module_inst_1_1845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5989]),.i2(intermediate_reg_0[5988]),.o(intermediate_reg_1[2994]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5987]),.i2(intermediate_reg_0[5986]),.o(intermediate_reg_1[2993]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5985]),.i2(intermediate_reg_0[5984]),.o(intermediate_reg_1[2992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5983]),.i2(intermediate_reg_0[5982]),.o(intermediate_reg_1[2991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5981]),.i2(intermediate_reg_0[5980]),.o(intermediate_reg_1[2990]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5979]),.i2(intermediate_reg_0[5978]),.o(intermediate_reg_1[2989]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5977]),.i2(intermediate_reg_0[5976]),.o(intermediate_reg_1[2988])); 
fsm fsm_inst_1_1852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5975]),.i2(intermediate_reg_0[5974]),.o(intermediate_reg_1[2987])); 
fsm fsm_inst_1_1853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5973]),.i2(intermediate_reg_0[5972]),.o(intermediate_reg_1[2986])); 
fsm fsm_inst_1_1854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5971]),.i2(intermediate_reg_0[5970]),.o(intermediate_reg_1[2985])); 
fsm fsm_inst_1_1855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5969]),.i2(intermediate_reg_0[5968]),.o(intermediate_reg_1[2984])); 
fsm fsm_inst_1_1856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5967]),.i2(intermediate_reg_0[5966]),.o(intermediate_reg_1[2983])); 
mux_module mux_module_inst_1_1857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5965]),.i2(intermediate_reg_0[5964]),.o(intermediate_reg_1[2982]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5963]),.i2(intermediate_reg_0[5962]),.o(intermediate_reg_1[2981])); 
fsm fsm_inst_1_1859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5961]),.i2(intermediate_reg_0[5960]),.o(intermediate_reg_1[2980])); 
fsm fsm_inst_1_1860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5959]),.i2(intermediate_reg_0[5958]),.o(intermediate_reg_1[2979])); 
fsm fsm_inst_1_1861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5957]),.i2(intermediate_reg_0[5956]),.o(intermediate_reg_1[2978])); 
fsm fsm_inst_1_1862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5955]),.i2(intermediate_reg_0[5954]),.o(intermediate_reg_1[2977])); 
mux_module mux_module_inst_1_1863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5953]),.i2(intermediate_reg_0[5952]),.o(intermediate_reg_1[2976]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5951]),.i2(intermediate_reg_0[5950]),.o(intermediate_reg_1[2975])); 
mux_module mux_module_inst_1_1865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5949]),.i2(intermediate_reg_0[5948]),.o(intermediate_reg_1[2974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5947]),.i2(intermediate_reg_0[5946]),.o(intermediate_reg_1[2973]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5945]),.i2(intermediate_reg_0[5944]),.o(intermediate_reg_1[2972])); 
fsm fsm_inst_1_1868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5943]),.i2(intermediate_reg_0[5942]),.o(intermediate_reg_1[2971])); 
mux_module mux_module_inst_1_1869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5941]),.i2(intermediate_reg_0[5940]),.o(intermediate_reg_1[2970]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5939]),.i2(intermediate_reg_0[5938]),.o(intermediate_reg_1[2969])); 
mux_module mux_module_inst_1_1871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5937]),.i2(intermediate_reg_0[5936]),.o(intermediate_reg_1[2968]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5935]),.i2(intermediate_reg_0[5934]),.o(intermediate_reg_1[2967])); 
fsm fsm_inst_1_1873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5933]),.i2(intermediate_reg_0[5932]),.o(intermediate_reg_1[2966])); 
fsm fsm_inst_1_1874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5931]),.i2(intermediate_reg_0[5930]),.o(intermediate_reg_1[2965])); 
mux_module mux_module_inst_1_1875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5929]),.i2(intermediate_reg_0[5928]),.o(intermediate_reg_1[2964]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5927]),.i2(intermediate_reg_0[5926]),.o(intermediate_reg_1[2963])); 
fsm fsm_inst_1_1877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5925]),.i2(intermediate_reg_0[5924]),.o(intermediate_reg_1[2962])); 
fsm fsm_inst_1_1878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5923]),.i2(intermediate_reg_0[5922]),.o(intermediate_reg_1[2961])); 
fsm fsm_inst_1_1879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5921]),.i2(intermediate_reg_0[5920]),.o(intermediate_reg_1[2960])); 
fsm fsm_inst_1_1880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5919]),.i2(intermediate_reg_0[5918]),.o(intermediate_reg_1[2959])); 
mux_module mux_module_inst_1_1881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5917]),.i2(intermediate_reg_0[5916]),.o(intermediate_reg_1[2958]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5915]),.i2(intermediate_reg_0[5914]),.o(intermediate_reg_1[2957])); 
fsm fsm_inst_1_1883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5913]),.i2(intermediate_reg_0[5912]),.o(intermediate_reg_1[2956])); 
mux_module mux_module_inst_1_1884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5911]),.i2(intermediate_reg_0[5910]),.o(intermediate_reg_1[2955]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5909]),.i2(intermediate_reg_0[5908]),.o(intermediate_reg_1[2954])); 
mux_module mux_module_inst_1_1886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5907]),.i2(intermediate_reg_0[5906]),.o(intermediate_reg_1[2953]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5905]),.i2(intermediate_reg_0[5904]),.o(intermediate_reg_1[2952]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5903]),.i2(intermediate_reg_0[5902]),.o(intermediate_reg_1[2951]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5901]),.i2(intermediate_reg_0[5900]),.o(intermediate_reg_1[2950])); 
fsm fsm_inst_1_1890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5899]),.i2(intermediate_reg_0[5898]),.o(intermediate_reg_1[2949])); 
fsm fsm_inst_1_1891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5897]),.i2(intermediate_reg_0[5896]),.o(intermediate_reg_1[2948])); 
fsm fsm_inst_1_1892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5895]),.i2(intermediate_reg_0[5894]),.o(intermediate_reg_1[2947])); 
fsm fsm_inst_1_1893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5893]),.i2(intermediate_reg_0[5892]),.o(intermediate_reg_1[2946])); 
fsm fsm_inst_1_1894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5891]),.i2(intermediate_reg_0[5890]),.o(intermediate_reg_1[2945])); 
fsm fsm_inst_1_1895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5889]),.i2(intermediate_reg_0[5888]),.o(intermediate_reg_1[2944])); 
mux_module mux_module_inst_1_1896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5887]),.i2(intermediate_reg_0[5886]),.o(intermediate_reg_1[2943]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5885]),.i2(intermediate_reg_0[5884]),.o(intermediate_reg_1[2942]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5883]),.i2(intermediate_reg_0[5882]),.o(intermediate_reg_1[2941])); 
mux_module mux_module_inst_1_1899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5881]),.i2(intermediate_reg_0[5880]),.o(intermediate_reg_1[2940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5879]),.i2(intermediate_reg_0[5878]),.o(intermediate_reg_1[2939]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5877]),.i2(intermediate_reg_0[5876]),.o(intermediate_reg_1[2938])); 
fsm fsm_inst_1_1902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5875]),.i2(intermediate_reg_0[5874]),.o(intermediate_reg_1[2937])); 
mux_module mux_module_inst_1_1903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5873]),.i2(intermediate_reg_0[5872]),.o(intermediate_reg_1[2936]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5871]),.i2(intermediate_reg_0[5870]),.o(intermediate_reg_1[2935])); 
mux_module mux_module_inst_1_1905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5869]),.i2(intermediate_reg_0[5868]),.o(intermediate_reg_1[2934]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5867]),.i2(intermediate_reg_0[5866]),.o(intermediate_reg_1[2933]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5865]),.i2(intermediate_reg_0[5864]),.o(intermediate_reg_1[2932]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5863]),.i2(intermediate_reg_0[5862]),.o(intermediate_reg_1[2931]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5861]),.i2(intermediate_reg_0[5860]),.o(intermediate_reg_1[2930])); 
mux_module mux_module_inst_1_1910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5859]),.i2(intermediate_reg_0[5858]),.o(intermediate_reg_1[2929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5857]),.i2(intermediate_reg_0[5856]),.o(intermediate_reg_1[2928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5855]),.i2(intermediate_reg_0[5854]),.o(intermediate_reg_1[2927]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5853]),.i2(intermediate_reg_0[5852]),.o(intermediate_reg_1[2926])); 
mux_module mux_module_inst_1_1914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5851]),.i2(intermediate_reg_0[5850]),.o(intermediate_reg_1[2925]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5849]),.i2(intermediate_reg_0[5848]),.o(intermediate_reg_1[2924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5847]),.i2(intermediate_reg_0[5846]),.o(intermediate_reg_1[2923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5845]),.i2(intermediate_reg_0[5844]),.o(intermediate_reg_1[2922]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5843]),.i2(intermediate_reg_0[5842]),.o(intermediate_reg_1[2921])); 
mux_module mux_module_inst_1_1919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5841]),.i2(intermediate_reg_0[5840]),.o(intermediate_reg_1[2920]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5839]),.i2(intermediate_reg_0[5838]),.o(intermediate_reg_1[2919])); 
mux_module mux_module_inst_1_1921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5837]),.i2(intermediate_reg_0[5836]),.o(intermediate_reg_1[2918]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5835]),.i2(intermediate_reg_0[5834]),.o(intermediate_reg_1[2917]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5833]),.i2(intermediate_reg_0[5832]),.o(intermediate_reg_1[2916])); 
mux_module mux_module_inst_1_1924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5831]),.i2(intermediate_reg_0[5830]),.o(intermediate_reg_1[2915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5829]),.i2(intermediate_reg_0[5828]),.o(intermediate_reg_1[2914]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5827]),.i2(intermediate_reg_0[5826]),.o(intermediate_reg_1[2913])); 
mux_module mux_module_inst_1_1927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5825]),.i2(intermediate_reg_0[5824]),.o(intermediate_reg_1[2912]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5823]),.i2(intermediate_reg_0[5822]),.o(intermediate_reg_1[2911]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5821]),.i2(intermediate_reg_0[5820]),.o(intermediate_reg_1[2910]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5819]),.i2(intermediate_reg_0[5818]),.o(intermediate_reg_1[2909]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5817]),.i2(intermediate_reg_0[5816]),.o(intermediate_reg_1[2908])); 
fsm fsm_inst_1_1932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5815]),.i2(intermediate_reg_0[5814]),.o(intermediate_reg_1[2907])); 
fsm fsm_inst_1_1933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5813]),.i2(intermediate_reg_0[5812]),.o(intermediate_reg_1[2906])); 
mux_module mux_module_inst_1_1934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5811]),.i2(intermediate_reg_0[5810]),.o(intermediate_reg_1[2905]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5809]),.i2(intermediate_reg_0[5808]),.o(intermediate_reg_1[2904])); 
fsm fsm_inst_1_1936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5807]),.i2(intermediate_reg_0[5806]),.o(intermediate_reg_1[2903])); 
fsm fsm_inst_1_1937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5805]),.i2(intermediate_reg_0[5804]),.o(intermediate_reg_1[2902])); 
mux_module mux_module_inst_1_1938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5803]),.i2(intermediate_reg_0[5802]),.o(intermediate_reg_1[2901]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5801]),.i2(intermediate_reg_0[5800]),.o(intermediate_reg_1[2900])); 
fsm fsm_inst_1_1940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5799]),.i2(intermediate_reg_0[5798]),.o(intermediate_reg_1[2899])); 
fsm fsm_inst_1_1941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5797]),.i2(intermediate_reg_0[5796]),.o(intermediate_reg_1[2898])); 
mux_module mux_module_inst_1_1942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5795]),.i2(intermediate_reg_0[5794]),.o(intermediate_reg_1[2897]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5793]),.i2(intermediate_reg_0[5792]),.o(intermediate_reg_1[2896])); 
fsm fsm_inst_1_1944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5791]),.i2(intermediate_reg_0[5790]),.o(intermediate_reg_1[2895])); 
mux_module mux_module_inst_1_1945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5789]),.i2(intermediate_reg_0[5788]),.o(intermediate_reg_1[2894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5787]),.i2(intermediate_reg_0[5786]),.o(intermediate_reg_1[2893]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5785]),.i2(intermediate_reg_0[5784]),.o(intermediate_reg_1[2892])); 
fsm fsm_inst_1_1948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5783]),.i2(intermediate_reg_0[5782]),.o(intermediate_reg_1[2891])); 
fsm fsm_inst_1_1949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5781]),.i2(intermediate_reg_0[5780]),.o(intermediate_reg_1[2890])); 
fsm fsm_inst_1_1950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5779]),.i2(intermediate_reg_0[5778]),.o(intermediate_reg_1[2889])); 
fsm fsm_inst_1_1951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5777]),.i2(intermediate_reg_0[5776]),.o(intermediate_reg_1[2888])); 
fsm fsm_inst_1_1952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5775]),.i2(intermediate_reg_0[5774]),.o(intermediate_reg_1[2887])); 
mux_module mux_module_inst_1_1953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5773]),.i2(intermediate_reg_0[5772]),.o(intermediate_reg_1[2886]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5771]),.i2(intermediate_reg_0[5770]),.o(intermediate_reg_1[2885]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5769]),.i2(intermediate_reg_0[5768]),.o(intermediate_reg_1[2884])); 
fsm fsm_inst_1_1956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5767]),.i2(intermediate_reg_0[5766]),.o(intermediate_reg_1[2883])); 
mux_module mux_module_inst_1_1957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5765]),.i2(intermediate_reg_0[5764]),.o(intermediate_reg_1[2882]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5763]),.i2(intermediate_reg_0[5762]),.o(intermediate_reg_1[2881]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5761]),.i2(intermediate_reg_0[5760]),.o(intermediate_reg_1[2880])); 
fsm fsm_inst_1_1960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5759]),.i2(intermediate_reg_0[5758]),.o(intermediate_reg_1[2879])); 
fsm fsm_inst_1_1961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5757]),.i2(intermediate_reg_0[5756]),.o(intermediate_reg_1[2878])); 
mux_module mux_module_inst_1_1962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5755]),.i2(intermediate_reg_0[5754]),.o(intermediate_reg_1[2877]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5753]),.i2(intermediate_reg_0[5752]),.o(intermediate_reg_1[2876]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5751]),.i2(intermediate_reg_0[5750]),.o(intermediate_reg_1[2875])); 
mux_module mux_module_inst_1_1965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5749]),.i2(intermediate_reg_0[5748]),.o(intermediate_reg_1[2874]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5747]),.i2(intermediate_reg_0[5746]),.o(intermediate_reg_1[2873])); 
mux_module mux_module_inst_1_1967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5745]),.i2(intermediate_reg_0[5744]),.o(intermediate_reg_1[2872]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5743]),.i2(intermediate_reg_0[5742]),.o(intermediate_reg_1[2871])); 
fsm fsm_inst_1_1969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5741]),.i2(intermediate_reg_0[5740]),.o(intermediate_reg_1[2870])); 
fsm fsm_inst_1_1970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5739]),.i2(intermediate_reg_0[5738]),.o(intermediate_reg_1[2869])); 
fsm fsm_inst_1_1971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5737]),.i2(intermediate_reg_0[5736]),.o(intermediate_reg_1[2868])); 
mux_module mux_module_inst_1_1972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5735]),.i2(intermediate_reg_0[5734]),.o(intermediate_reg_1[2867]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5733]),.i2(intermediate_reg_0[5732]),.o(intermediate_reg_1[2866])); 
fsm fsm_inst_1_1974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5731]),.i2(intermediate_reg_0[5730]),.o(intermediate_reg_1[2865])); 
mux_module mux_module_inst_1_1975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5729]),.i2(intermediate_reg_0[5728]),.o(intermediate_reg_1[2864]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5727]),.i2(intermediate_reg_0[5726]),.o(intermediate_reg_1[2863]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5725]),.i2(intermediate_reg_0[5724]),.o(intermediate_reg_1[2862]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5723]),.i2(intermediate_reg_0[5722]),.o(intermediate_reg_1[2861])); 
mux_module mux_module_inst_1_1979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5721]),.i2(intermediate_reg_0[5720]),.o(intermediate_reg_1[2860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5719]),.i2(intermediate_reg_0[5718]),.o(intermediate_reg_1[2859]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5717]),.i2(intermediate_reg_0[5716]),.o(intermediate_reg_1[2858])); 
fsm fsm_inst_1_1982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5715]),.i2(intermediate_reg_0[5714]),.o(intermediate_reg_1[2857])); 
mux_module mux_module_inst_1_1983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5713]),.i2(intermediate_reg_0[5712]),.o(intermediate_reg_1[2856]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5711]),.i2(intermediate_reg_0[5710]),.o(intermediate_reg_1[2855])); 
fsm fsm_inst_1_1985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5709]),.i2(intermediate_reg_0[5708]),.o(intermediate_reg_1[2854])); 
fsm fsm_inst_1_1986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5707]),.i2(intermediate_reg_0[5706]),.o(intermediate_reg_1[2853])); 
fsm fsm_inst_1_1987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5705]),.i2(intermediate_reg_0[5704]),.o(intermediate_reg_1[2852])); 
mux_module mux_module_inst_1_1988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5703]),.i2(intermediate_reg_0[5702]),.o(intermediate_reg_1[2851]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5701]),.i2(intermediate_reg_0[5700]),.o(intermediate_reg_1[2850])); 
mux_module mux_module_inst_1_1990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5699]),.i2(intermediate_reg_0[5698]),.o(intermediate_reg_1[2849]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5697]),.i2(intermediate_reg_0[5696]),.o(intermediate_reg_1[2848])); 
fsm fsm_inst_1_1992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5695]),.i2(intermediate_reg_0[5694]),.o(intermediate_reg_1[2847])); 
fsm fsm_inst_1_1993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5693]),.i2(intermediate_reg_0[5692]),.o(intermediate_reg_1[2846])); 
fsm fsm_inst_1_1994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5691]),.i2(intermediate_reg_0[5690]),.o(intermediate_reg_1[2845])); 
fsm fsm_inst_1_1995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5689]),.i2(intermediate_reg_0[5688]),.o(intermediate_reg_1[2844])); 
mux_module mux_module_inst_1_1996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5687]),.i2(intermediate_reg_0[5686]),.o(intermediate_reg_1[2843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5685]),.i2(intermediate_reg_0[5684]),.o(intermediate_reg_1[2842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5683]),.i2(intermediate_reg_0[5682]),.o(intermediate_reg_1[2841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5681]),.i2(intermediate_reg_0[5680]),.o(intermediate_reg_1[2840]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5679]),.i2(intermediate_reg_0[5678]),.o(intermediate_reg_1[2839]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5677]),.i2(intermediate_reg_0[5676]),.o(intermediate_reg_1[2838])); 
fsm fsm_inst_1_2002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5675]),.i2(intermediate_reg_0[5674]),.o(intermediate_reg_1[2837])); 
mux_module mux_module_inst_1_2003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5673]),.i2(intermediate_reg_0[5672]),.o(intermediate_reg_1[2836]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5671]),.i2(intermediate_reg_0[5670]),.o(intermediate_reg_1[2835])); 
mux_module mux_module_inst_1_2005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5669]),.i2(intermediate_reg_0[5668]),.o(intermediate_reg_1[2834]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5667]),.i2(intermediate_reg_0[5666]),.o(intermediate_reg_1[2833]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5665]),.i2(intermediate_reg_0[5664]),.o(intermediate_reg_1[2832]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5663]),.i2(intermediate_reg_0[5662]),.o(intermediate_reg_1[2831]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5661]),.i2(intermediate_reg_0[5660]),.o(intermediate_reg_1[2830])); 
mux_module mux_module_inst_1_2010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5659]),.i2(intermediate_reg_0[5658]),.o(intermediate_reg_1[2829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5657]),.i2(intermediate_reg_0[5656]),.o(intermediate_reg_1[2828]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5655]),.i2(intermediate_reg_0[5654]),.o(intermediate_reg_1[2827]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5653]),.i2(intermediate_reg_0[5652]),.o(intermediate_reg_1[2826]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5651]),.i2(intermediate_reg_0[5650]),.o(intermediate_reg_1[2825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5649]),.i2(intermediate_reg_0[5648]),.o(intermediate_reg_1[2824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5647]),.i2(intermediate_reg_0[5646]),.o(intermediate_reg_1[2823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5645]),.i2(intermediate_reg_0[5644]),.o(intermediate_reg_1[2822]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5643]),.i2(intermediate_reg_0[5642]),.o(intermediate_reg_1[2821]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5641]),.i2(intermediate_reg_0[5640]),.o(intermediate_reg_1[2820])); 
fsm fsm_inst_1_2020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5639]),.i2(intermediate_reg_0[5638]),.o(intermediate_reg_1[2819])); 
mux_module mux_module_inst_1_2021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5637]),.i2(intermediate_reg_0[5636]),.o(intermediate_reg_1[2818]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5635]),.i2(intermediate_reg_0[5634]),.o(intermediate_reg_1[2817])); 
mux_module mux_module_inst_1_2023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5633]),.i2(intermediate_reg_0[5632]),.o(intermediate_reg_1[2816]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5631]),.i2(intermediate_reg_0[5630]),.o(intermediate_reg_1[2815]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5629]),.i2(intermediate_reg_0[5628]),.o(intermediate_reg_1[2814])); 
fsm fsm_inst_1_2026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5627]),.i2(intermediate_reg_0[5626]),.o(intermediate_reg_1[2813])); 
fsm fsm_inst_1_2027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5625]),.i2(intermediate_reg_0[5624]),.o(intermediate_reg_1[2812])); 
mux_module mux_module_inst_1_2028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5623]),.i2(intermediate_reg_0[5622]),.o(intermediate_reg_1[2811]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5621]),.i2(intermediate_reg_0[5620]),.o(intermediate_reg_1[2810])); 
fsm fsm_inst_1_2030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5619]),.i2(intermediate_reg_0[5618]),.o(intermediate_reg_1[2809])); 
fsm fsm_inst_1_2031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5617]),.i2(intermediate_reg_0[5616]),.o(intermediate_reg_1[2808])); 
fsm fsm_inst_1_2032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5615]),.i2(intermediate_reg_0[5614]),.o(intermediate_reg_1[2807])); 
fsm fsm_inst_1_2033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5613]),.i2(intermediate_reg_0[5612]),.o(intermediate_reg_1[2806])); 
fsm fsm_inst_1_2034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5611]),.i2(intermediate_reg_0[5610]),.o(intermediate_reg_1[2805])); 
mux_module mux_module_inst_1_2035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5609]),.i2(intermediate_reg_0[5608]),.o(intermediate_reg_1[2804]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5607]),.i2(intermediate_reg_0[5606]),.o(intermediate_reg_1[2803])); 
mux_module mux_module_inst_1_2037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5605]),.i2(intermediate_reg_0[5604]),.o(intermediate_reg_1[2802]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5603]),.i2(intermediate_reg_0[5602]),.o(intermediate_reg_1[2801]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5601]),.i2(intermediate_reg_0[5600]),.o(intermediate_reg_1[2800])); 
mux_module mux_module_inst_1_2040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5599]),.i2(intermediate_reg_0[5598]),.o(intermediate_reg_1[2799]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5597]),.i2(intermediate_reg_0[5596]),.o(intermediate_reg_1[2798]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5595]),.i2(intermediate_reg_0[5594]),.o(intermediate_reg_1[2797]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5593]),.i2(intermediate_reg_0[5592]),.o(intermediate_reg_1[2796])); 
mux_module mux_module_inst_1_2044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5591]),.i2(intermediate_reg_0[5590]),.o(intermediate_reg_1[2795]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5589]),.i2(intermediate_reg_0[5588]),.o(intermediate_reg_1[2794])); 
mux_module mux_module_inst_1_2046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5587]),.i2(intermediate_reg_0[5586]),.o(intermediate_reg_1[2793]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5585]),.i2(intermediate_reg_0[5584]),.o(intermediate_reg_1[2792]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5583]),.i2(intermediate_reg_0[5582]),.o(intermediate_reg_1[2791]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5581]),.i2(intermediate_reg_0[5580]),.o(intermediate_reg_1[2790]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5579]),.i2(intermediate_reg_0[5578]),.o(intermediate_reg_1[2789]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5577]),.i2(intermediate_reg_0[5576]),.o(intermediate_reg_1[2788])); 
mux_module mux_module_inst_1_2052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5575]),.i2(intermediate_reg_0[5574]),.o(intermediate_reg_1[2787]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5573]),.i2(intermediate_reg_0[5572]),.o(intermediate_reg_1[2786]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5571]),.i2(intermediate_reg_0[5570]),.o(intermediate_reg_1[2785])); 
mux_module mux_module_inst_1_2055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5569]),.i2(intermediate_reg_0[5568]),.o(intermediate_reg_1[2784]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5567]),.i2(intermediate_reg_0[5566]),.o(intermediate_reg_1[2783]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5565]),.i2(intermediate_reg_0[5564]),.o(intermediate_reg_1[2782])); 
mux_module mux_module_inst_1_2058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5563]),.i2(intermediate_reg_0[5562]),.o(intermediate_reg_1[2781]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5561]),.i2(intermediate_reg_0[5560]),.o(intermediate_reg_1[2780])); 
mux_module mux_module_inst_1_2060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5559]),.i2(intermediate_reg_0[5558]),.o(intermediate_reg_1[2779]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5557]),.i2(intermediate_reg_0[5556]),.o(intermediate_reg_1[2778]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5555]),.i2(intermediate_reg_0[5554]),.o(intermediate_reg_1[2777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5553]),.i2(intermediate_reg_0[5552]),.o(intermediate_reg_1[2776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5551]),.i2(intermediate_reg_0[5550]),.o(intermediate_reg_1[2775]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5549]),.i2(intermediate_reg_0[5548]),.o(intermediate_reg_1[2774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5547]),.i2(intermediate_reg_0[5546]),.o(intermediate_reg_1[2773]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5545]),.i2(intermediate_reg_0[5544]),.o(intermediate_reg_1[2772])); 
fsm fsm_inst_1_2068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5543]),.i2(intermediate_reg_0[5542]),.o(intermediate_reg_1[2771])); 
mux_module mux_module_inst_1_2069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5541]),.i2(intermediate_reg_0[5540]),.o(intermediate_reg_1[2770]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5539]),.i2(intermediate_reg_0[5538]),.o(intermediate_reg_1[2769])); 
mux_module mux_module_inst_1_2071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5537]),.i2(intermediate_reg_0[5536]),.o(intermediate_reg_1[2768]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5535]),.i2(intermediate_reg_0[5534]),.o(intermediate_reg_1[2767])); 
fsm fsm_inst_1_2073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5533]),.i2(intermediate_reg_0[5532]),.o(intermediate_reg_1[2766])); 
mux_module mux_module_inst_1_2074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5531]),.i2(intermediate_reg_0[5530]),.o(intermediate_reg_1[2765]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5529]),.i2(intermediate_reg_0[5528]),.o(intermediate_reg_1[2764])); 
fsm fsm_inst_1_2076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5527]),.i2(intermediate_reg_0[5526]),.o(intermediate_reg_1[2763])); 
mux_module mux_module_inst_1_2077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5525]),.i2(intermediate_reg_0[5524]),.o(intermediate_reg_1[2762]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5523]),.i2(intermediate_reg_0[5522]),.o(intermediate_reg_1[2761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5521]),.i2(intermediate_reg_0[5520]),.o(intermediate_reg_1[2760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5519]),.i2(intermediate_reg_0[5518]),.o(intermediate_reg_1[2759]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5517]),.i2(intermediate_reg_0[5516]),.o(intermediate_reg_1[2758])); 
fsm fsm_inst_1_2082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5515]),.i2(intermediate_reg_0[5514]),.o(intermediate_reg_1[2757])); 
fsm fsm_inst_1_2083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5513]),.i2(intermediate_reg_0[5512]),.o(intermediate_reg_1[2756])); 
mux_module mux_module_inst_1_2084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5511]),.i2(intermediate_reg_0[5510]),.o(intermediate_reg_1[2755]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5509]),.i2(intermediate_reg_0[5508]),.o(intermediate_reg_1[2754])); 
fsm fsm_inst_1_2086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5507]),.i2(intermediate_reg_0[5506]),.o(intermediate_reg_1[2753])); 
fsm fsm_inst_1_2087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5505]),.i2(intermediate_reg_0[5504]),.o(intermediate_reg_1[2752])); 
mux_module mux_module_inst_1_2088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5503]),.i2(intermediate_reg_0[5502]),.o(intermediate_reg_1[2751]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5501]),.i2(intermediate_reg_0[5500]),.o(intermediate_reg_1[2750])); 
mux_module mux_module_inst_1_2090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5499]),.i2(intermediate_reg_0[5498]),.o(intermediate_reg_1[2749]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5497]),.i2(intermediate_reg_0[5496]),.o(intermediate_reg_1[2748])); 
fsm fsm_inst_1_2092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5495]),.i2(intermediate_reg_0[5494]),.o(intermediate_reg_1[2747])); 
mux_module mux_module_inst_1_2093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5493]),.i2(intermediate_reg_0[5492]),.o(intermediate_reg_1[2746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5491]),.i2(intermediate_reg_0[5490]),.o(intermediate_reg_1[2745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5489]),.i2(intermediate_reg_0[5488]),.o(intermediate_reg_1[2744]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5487]),.i2(intermediate_reg_0[5486]),.o(intermediate_reg_1[2743])); 
mux_module mux_module_inst_1_2097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5485]),.i2(intermediate_reg_0[5484]),.o(intermediate_reg_1[2742]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5483]),.i2(intermediate_reg_0[5482]),.o(intermediate_reg_1[2741])); 
fsm fsm_inst_1_2099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5481]),.i2(intermediate_reg_0[5480]),.o(intermediate_reg_1[2740])); 
mux_module mux_module_inst_1_2100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5479]),.i2(intermediate_reg_0[5478]),.o(intermediate_reg_1[2739]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5477]),.i2(intermediate_reg_0[5476]),.o(intermediate_reg_1[2738])); 
fsm fsm_inst_1_2102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5475]),.i2(intermediate_reg_0[5474]),.o(intermediate_reg_1[2737])); 
mux_module mux_module_inst_1_2103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5473]),.i2(intermediate_reg_0[5472]),.o(intermediate_reg_1[2736]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5471]),.i2(intermediate_reg_0[5470]),.o(intermediate_reg_1[2735]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5469]),.i2(intermediate_reg_0[5468]),.o(intermediate_reg_1[2734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5467]),.i2(intermediate_reg_0[5466]),.o(intermediate_reg_1[2733]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5465]),.i2(intermediate_reg_0[5464]),.o(intermediate_reg_1[2732]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5463]),.i2(intermediate_reg_0[5462]),.o(intermediate_reg_1[2731])); 
mux_module mux_module_inst_1_2109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5461]),.i2(intermediate_reg_0[5460]),.o(intermediate_reg_1[2730]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5459]),.i2(intermediate_reg_0[5458]),.o(intermediate_reg_1[2729])); 
fsm fsm_inst_1_2111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5457]),.i2(intermediate_reg_0[5456]),.o(intermediate_reg_1[2728])); 
mux_module mux_module_inst_1_2112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5455]),.i2(intermediate_reg_0[5454]),.o(intermediate_reg_1[2727]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5453]),.i2(intermediate_reg_0[5452]),.o(intermediate_reg_1[2726])); 
fsm fsm_inst_1_2114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5451]),.i2(intermediate_reg_0[5450]),.o(intermediate_reg_1[2725])); 
fsm fsm_inst_1_2115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5449]),.i2(intermediate_reg_0[5448]),.o(intermediate_reg_1[2724])); 
mux_module mux_module_inst_1_2116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5447]),.i2(intermediate_reg_0[5446]),.o(intermediate_reg_1[2723]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5445]),.i2(intermediate_reg_0[5444]),.o(intermediate_reg_1[2722]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5443]),.i2(intermediate_reg_0[5442]),.o(intermediate_reg_1[2721]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5441]),.i2(intermediate_reg_0[5440]),.o(intermediate_reg_1[2720])); 
fsm fsm_inst_1_2120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5439]),.i2(intermediate_reg_0[5438]),.o(intermediate_reg_1[2719])); 
mux_module mux_module_inst_1_2121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5437]),.i2(intermediate_reg_0[5436]),.o(intermediate_reg_1[2718]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5435]),.i2(intermediate_reg_0[5434]),.o(intermediate_reg_1[2717])); 
fsm fsm_inst_1_2123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5433]),.i2(intermediate_reg_0[5432]),.o(intermediate_reg_1[2716])); 
mux_module mux_module_inst_1_2124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5431]),.i2(intermediate_reg_0[5430]),.o(intermediate_reg_1[2715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5429]),.i2(intermediate_reg_0[5428]),.o(intermediate_reg_1[2714]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5427]),.i2(intermediate_reg_0[5426]),.o(intermediate_reg_1[2713]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5425]),.i2(intermediate_reg_0[5424]),.o(intermediate_reg_1[2712])); 
fsm fsm_inst_1_2128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5423]),.i2(intermediate_reg_0[5422]),.o(intermediate_reg_1[2711])); 
mux_module mux_module_inst_1_2129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5421]),.i2(intermediate_reg_0[5420]),.o(intermediate_reg_1[2710]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5419]),.i2(intermediate_reg_0[5418]),.o(intermediate_reg_1[2709])); 
fsm fsm_inst_1_2131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5417]),.i2(intermediate_reg_0[5416]),.o(intermediate_reg_1[2708])); 
fsm fsm_inst_1_2132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5415]),.i2(intermediate_reg_0[5414]),.o(intermediate_reg_1[2707])); 
mux_module mux_module_inst_1_2133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5413]),.i2(intermediate_reg_0[5412]),.o(intermediate_reg_1[2706]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5411]),.i2(intermediate_reg_0[5410]),.o(intermediate_reg_1[2705])); 
fsm fsm_inst_1_2135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5409]),.i2(intermediate_reg_0[5408]),.o(intermediate_reg_1[2704])); 
fsm fsm_inst_1_2136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5407]),.i2(intermediate_reg_0[5406]),.o(intermediate_reg_1[2703])); 
mux_module mux_module_inst_1_2137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5405]),.i2(intermediate_reg_0[5404]),.o(intermediate_reg_1[2702]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5403]),.i2(intermediate_reg_0[5402]),.o(intermediate_reg_1[2701]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5401]),.i2(intermediate_reg_0[5400]),.o(intermediate_reg_1[2700])); 
mux_module mux_module_inst_1_2140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5399]),.i2(intermediate_reg_0[5398]),.o(intermediate_reg_1[2699]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5397]),.i2(intermediate_reg_0[5396]),.o(intermediate_reg_1[2698])); 
mux_module mux_module_inst_1_2142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5395]),.i2(intermediate_reg_0[5394]),.o(intermediate_reg_1[2697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5393]),.i2(intermediate_reg_0[5392]),.o(intermediate_reg_1[2696]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5391]),.i2(intermediate_reg_0[5390]),.o(intermediate_reg_1[2695]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5389]),.i2(intermediate_reg_0[5388]),.o(intermediate_reg_1[2694]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5387]),.i2(intermediate_reg_0[5386]),.o(intermediate_reg_1[2693])); 
fsm fsm_inst_1_2147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5385]),.i2(intermediate_reg_0[5384]),.o(intermediate_reg_1[2692])); 
fsm fsm_inst_1_2148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5383]),.i2(intermediate_reg_0[5382]),.o(intermediate_reg_1[2691])); 
fsm fsm_inst_1_2149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5381]),.i2(intermediate_reg_0[5380]),.o(intermediate_reg_1[2690])); 
mux_module mux_module_inst_1_2150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5379]),.i2(intermediate_reg_0[5378]),.o(intermediate_reg_1[2689]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5377]),.i2(intermediate_reg_0[5376]),.o(intermediate_reg_1[2688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5375]),.i2(intermediate_reg_0[5374]),.o(intermediate_reg_1[2687]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5373]),.i2(intermediate_reg_0[5372]),.o(intermediate_reg_1[2686])); 
fsm fsm_inst_1_2154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5371]),.i2(intermediate_reg_0[5370]),.o(intermediate_reg_1[2685])); 
mux_module mux_module_inst_1_2155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5369]),.i2(intermediate_reg_0[5368]),.o(intermediate_reg_1[2684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5367]),.i2(intermediate_reg_0[5366]),.o(intermediate_reg_1[2683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5365]),.i2(intermediate_reg_0[5364]),.o(intermediate_reg_1[2682]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5363]),.i2(intermediate_reg_0[5362]),.o(intermediate_reg_1[2681])); 
mux_module mux_module_inst_1_2159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5361]),.i2(intermediate_reg_0[5360]),.o(intermediate_reg_1[2680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5359]),.i2(intermediate_reg_0[5358]),.o(intermediate_reg_1[2679]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5357]),.i2(intermediate_reg_0[5356]),.o(intermediate_reg_1[2678]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5355]),.i2(intermediate_reg_0[5354]),.o(intermediate_reg_1[2677])); 
mux_module mux_module_inst_1_2163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5353]),.i2(intermediate_reg_0[5352]),.o(intermediate_reg_1[2676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5351]),.i2(intermediate_reg_0[5350]),.o(intermediate_reg_1[2675]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5349]),.i2(intermediate_reg_0[5348]),.o(intermediate_reg_1[2674])); 
mux_module mux_module_inst_1_2166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5347]),.i2(intermediate_reg_0[5346]),.o(intermediate_reg_1[2673]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5345]),.i2(intermediate_reg_0[5344]),.o(intermediate_reg_1[2672]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5343]),.i2(intermediate_reg_0[5342]),.o(intermediate_reg_1[2671])); 
mux_module mux_module_inst_1_2169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5341]),.i2(intermediate_reg_0[5340]),.o(intermediate_reg_1[2670]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5339]),.i2(intermediate_reg_0[5338]),.o(intermediate_reg_1[2669]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5337]),.i2(intermediate_reg_0[5336]),.o(intermediate_reg_1[2668]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5335]),.i2(intermediate_reg_0[5334]),.o(intermediate_reg_1[2667])); 
fsm fsm_inst_1_2173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5333]),.i2(intermediate_reg_0[5332]),.o(intermediate_reg_1[2666])); 
mux_module mux_module_inst_1_2174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5331]),.i2(intermediate_reg_0[5330]),.o(intermediate_reg_1[2665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5329]),.i2(intermediate_reg_0[5328]),.o(intermediate_reg_1[2664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5327]),.i2(intermediate_reg_0[5326]),.o(intermediate_reg_1[2663]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5325]),.i2(intermediate_reg_0[5324]),.o(intermediate_reg_1[2662]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5323]),.i2(intermediate_reg_0[5322]),.o(intermediate_reg_1[2661])); 
mux_module mux_module_inst_1_2179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5321]),.i2(intermediate_reg_0[5320]),.o(intermediate_reg_1[2660]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5319]),.i2(intermediate_reg_0[5318]),.o(intermediate_reg_1[2659])); 
fsm fsm_inst_1_2181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5317]),.i2(intermediate_reg_0[5316]),.o(intermediate_reg_1[2658])); 
fsm fsm_inst_1_2182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5315]),.i2(intermediate_reg_0[5314]),.o(intermediate_reg_1[2657])); 
fsm fsm_inst_1_2183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5313]),.i2(intermediate_reg_0[5312]),.o(intermediate_reg_1[2656])); 
fsm fsm_inst_1_2184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5311]),.i2(intermediate_reg_0[5310]),.o(intermediate_reg_1[2655])); 
fsm fsm_inst_1_2185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5309]),.i2(intermediate_reg_0[5308]),.o(intermediate_reg_1[2654])); 
fsm fsm_inst_1_2186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5307]),.i2(intermediate_reg_0[5306]),.o(intermediate_reg_1[2653])); 
fsm fsm_inst_1_2187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5305]),.i2(intermediate_reg_0[5304]),.o(intermediate_reg_1[2652])); 
fsm fsm_inst_1_2188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5303]),.i2(intermediate_reg_0[5302]),.o(intermediate_reg_1[2651])); 
mux_module mux_module_inst_1_2189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5301]),.i2(intermediate_reg_0[5300]),.o(intermediate_reg_1[2650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5299]),.i2(intermediate_reg_0[5298]),.o(intermediate_reg_1[2649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5297]),.i2(intermediate_reg_0[5296]),.o(intermediate_reg_1[2648]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5295]),.i2(intermediate_reg_0[5294]),.o(intermediate_reg_1[2647])); 
mux_module mux_module_inst_1_2193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5293]),.i2(intermediate_reg_0[5292]),.o(intermediate_reg_1[2646]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5291]),.i2(intermediate_reg_0[5290]),.o(intermediate_reg_1[2645])); 
mux_module mux_module_inst_1_2195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5289]),.i2(intermediate_reg_0[5288]),.o(intermediate_reg_1[2644]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5287]),.i2(intermediate_reg_0[5286]),.o(intermediate_reg_1[2643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5285]),.i2(intermediate_reg_0[5284]),.o(intermediate_reg_1[2642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5283]),.i2(intermediate_reg_0[5282]),.o(intermediate_reg_1[2641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5281]),.i2(intermediate_reg_0[5280]),.o(intermediate_reg_1[2640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5279]),.i2(intermediate_reg_0[5278]),.o(intermediate_reg_1[2639]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5277]),.i2(intermediate_reg_0[5276]),.o(intermediate_reg_1[2638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5275]),.i2(intermediate_reg_0[5274]),.o(intermediate_reg_1[2637])); 
fsm fsm_inst_1_2203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5273]),.i2(intermediate_reg_0[5272]),.o(intermediate_reg_1[2636])); 
fsm fsm_inst_1_2204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5271]),.i2(intermediate_reg_0[5270]),.o(intermediate_reg_1[2635])); 
fsm fsm_inst_1_2205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5269]),.i2(intermediate_reg_0[5268]),.o(intermediate_reg_1[2634])); 
mux_module mux_module_inst_1_2206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5267]),.i2(intermediate_reg_0[5266]),.o(intermediate_reg_1[2633]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5265]),.i2(intermediate_reg_0[5264]),.o(intermediate_reg_1[2632])); 
mux_module mux_module_inst_1_2208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5263]),.i2(intermediate_reg_0[5262]),.o(intermediate_reg_1[2631]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5261]),.i2(intermediate_reg_0[5260]),.o(intermediate_reg_1[2630])); 
fsm fsm_inst_1_2210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5259]),.i2(intermediate_reg_0[5258]),.o(intermediate_reg_1[2629])); 
mux_module mux_module_inst_1_2211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5257]),.i2(intermediate_reg_0[5256]),.o(intermediate_reg_1[2628]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5255]),.i2(intermediate_reg_0[5254]),.o(intermediate_reg_1[2627])); 
mux_module mux_module_inst_1_2213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5253]),.i2(intermediate_reg_0[5252]),.o(intermediate_reg_1[2626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5251]),.i2(intermediate_reg_0[5250]),.o(intermediate_reg_1[2625])); 
fsm fsm_inst_1_2215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5249]),.i2(intermediate_reg_0[5248]),.o(intermediate_reg_1[2624])); 
mux_module mux_module_inst_1_2216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5247]),.i2(intermediate_reg_0[5246]),.o(intermediate_reg_1[2623]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5245]),.i2(intermediate_reg_0[5244]),.o(intermediate_reg_1[2622]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5243]),.i2(intermediate_reg_0[5242]),.o(intermediate_reg_1[2621])); 
fsm fsm_inst_1_2219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5241]),.i2(intermediate_reg_0[5240]),.o(intermediate_reg_1[2620])); 
fsm fsm_inst_1_2220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5239]),.i2(intermediate_reg_0[5238]),.o(intermediate_reg_1[2619])); 
fsm fsm_inst_1_2221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5237]),.i2(intermediate_reg_0[5236]),.o(intermediate_reg_1[2618])); 
fsm fsm_inst_1_2222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5235]),.i2(intermediate_reg_0[5234]),.o(intermediate_reg_1[2617])); 
mux_module mux_module_inst_1_2223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5233]),.i2(intermediate_reg_0[5232]),.o(intermediate_reg_1[2616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5231]),.i2(intermediate_reg_0[5230]),.o(intermediate_reg_1[2615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5229]),.i2(intermediate_reg_0[5228]),.o(intermediate_reg_1[2614]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5227]),.i2(intermediate_reg_0[5226]),.o(intermediate_reg_1[2613])); 
fsm fsm_inst_1_2227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5225]),.i2(intermediate_reg_0[5224]),.o(intermediate_reg_1[2612])); 
mux_module mux_module_inst_1_2228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5223]),.i2(intermediate_reg_0[5222]),.o(intermediate_reg_1[2611]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5221]),.i2(intermediate_reg_0[5220]),.o(intermediate_reg_1[2610])); 
mux_module mux_module_inst_1_2230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5219]),.i2(intermediate_reg_0[5218]),.o(intermediate_reg_1[2609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5217]),.i2(intermediate_reg_0[5216]),.o(intermediate_reg_1[2608]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5215]),.i2(intermediate_reg_0[5214]),.o(intermediate_reg_1[2607])); 
mux_module mux_module_inst_1_2233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5213]),.i2(intermediate_reg_0[5212]),.o(intermediate_reg_1[2606]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5211]),.i2(intermediate_reg_0[5210]),.o(intermediate_reg_1[2605])); 
fsm fsm_inst_1_2235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5209]),.i2(intermediate_reg_0[5208]),.o(intermediate_reg_1[2604])); 
fsm fsm_inst_1_2236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5207]),.i2(intermediate_reg_0[5206]),.o(intermediate_reg_1[2603])); 
mux_module mux_module_inst_1_2237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5205]),.i2(intermediate_reg_0[5204]),.o(intermediate_reg_1[2602]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5203]),.i2(intermediate_reg_0[5202]),.o(intermediate_reg_1[2601]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5201]),.i2(intermediate_reg_0[5200]),.o(intermediate_reg_1[2600]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5199]),.i2(intermediate_reg_0[5198]),.o(intermediate_reg_1[2599]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5197]),.i2(intermediate_reg_0[5196]),.o(intermediate_reg_1[2598]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5195]),.i2(intermediate_reg_0[5194]),.o(intermediate_reg_1[2597])); 
mux_module mux_module_inst_1_2243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5193]),.i2(intermediate_reg_0[5192]),.o(intermediate_reg_1[2596]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5191]),.i2(intermediate_reg_0[5190]),.o(intermediate_reg_1[2595])); 
fsm fsm_inst_1_2245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5189]),.i2(intermediate_reg_0[5188]),.o(intermediate_reg_1[2594])); 
fsm fsm_inst_1_2246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5187]),.i2(intermediate_reg_0[5186]),.o(intermediate_reg_1[2593])); 
mux_module mux_module_inst_1_2247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5185]),.i2(intermediate_reg_0[5184]),.o(intermediate_reg_1[2592]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5183]),.i2(intermediate_reg_0[5182]),.o(intermediate_reg_1[2591])); 
fsm fsm_inst_1_2249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5181]),.i2(intermediate_reg_0[5180]),.o(intermediate_reg_1[2590])); 
fsm fsm_inst_1_2250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5179]),.i2(intermediate_reg_0[5178]),.o(intermediate_reg_1[2589])); 
mux_module mux_module_inst_1_2251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5177]),.i2(intermediate_reg_0[5176]),.o(intermediate_reg_1[2588]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5175]),.i2(intermediate_reg_0[5174]),.o(intermediate_reg_1[2587])); 
fsm fsm_inst_1_2253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5173]),.i2(intermediate_reg_0[5172]),.o(intermediate_reg_1[2586])); 
fsm fsm_inst_1_2254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5171]),.i2(intermediate_reg_0[5170]),.o(intermediate_reg_1[2585])); 
fsm fsm_inst_1_2255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5169]),.i2(intermediate_reg_0[5168]),.o(intermediate_reg_1[2584])); 
fsm fsm_inst_1_2256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5167]),.i2(intermediate_reg_0[5166]),.o(intermediate_reg_1[2583])); 
fsm fsm_inst_1_2257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5165]),.i2(intermediate_reg_0[5164]),.o(intermediate_reg_1[2582])); 
mux_module mux_module_inst_1_2258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5163]),.i2(intermediate_reg_0[5162]),.o(intermediate_reg_1[2581]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5161]),.i2(intermediate_reg_0[5160]),.o(intermediate_reg_1[2580]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5159]),.i2(intermediate_reg_0[5158]),.o(intermediate_reg_1[2579]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5157]),.i2(intermediate_reg_0[5156]),.o(intermediate_reg_1[2578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5155]),.i2(intermediate_reg_0[5154]),.o(intermediate_reg_1[2577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5153]),.i2(intermediate_reg_0[5152]),.o(intermediate_reg_1[2576]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5151]),.i2(intermediate_reg_0[5150]),.o(intermediate_reg_1[2575]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5149]),.i2(intermediate_reg_0[5148]),.o(intermediate_reg_1[2574])); 
fsm fsm_inst_1_2266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5147]),.i2(intermediate_reg_0[5146]),.o(intermediate_reg_1[2573])); 
mux_module mux_module_inst_1_2267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5145]),.i2(intermediate_reg_0[5144]),.o(intermediate_reg_1[2572]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5143]),.i2(intermediate_reg_0[5142]),.o(intermediate_reg_1[2571])); 
fsm fsm_inst_1_2269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5141]),.i2(intermediate_reg_0[5140]),.o(intermediate_reg_1[2570])); 
mux_module mux_module_inst_1_2270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5139]),.i2(intermediate_reg_0[5138]),.o(intermediate_reg_1[2569]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5137]),.i2(intermediate_reg_0[5136]),.o(intermediate_reg_1[2568])); 
fsm fsm_inst_1_2272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5135]),.i2(intermediate_reg_0[5134]),.o(intermediate_reg_1[2567])); 
fsm fsm_inst_1_2273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5133]),.i2(intermediate_reg_0[5132]),.o(intermediate_reg_1[2566])); 
fsm fsm_inst_1_2274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5131]),.i2(intermediate_reg_0[5130]),.o(intermediate_reg_1[2565])); 
fsm fsm_inst_1_2275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5129]),.i2(intermediate_reg_0[5128]),.o(intermediate_reg_1[2564])); 
fsm fsm_inst_1_2276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5127]),.i2(intermediate_reg_0[5126]),.o(intermediate_reg_1[2563])); 
fsm fsm_inst_1_2277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5125]),.i2(intermediate_reg_0[5124]),.o(intermediate_reg_1[2562])); 
fsm fsm_inst_1_2278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5123]),.i2(intermediate_reg_0[5122]),.o(intermediate_reg_1[2561])); 
mux_module mux_module_inst_1_2279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5121]),.i2(intermediate_reg_0[5120]),.o(intermediate_reg_1[2560]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5119]),.i2(intermediate_reg_0[5118]),.o(intermediate_reg_1[2559]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5117]),.i2(intermediate_reg_0[5116]),.o(intermediate_reg_1[2558])); 
mux_module mux_module_inst_1_2282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5115]),.i2(intermediate_reg_0[5114]),.o(intermediate_reg_1[2557]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5113]),.i2(intermediate_reg_0[5112]),.o(intermediate_reg_1[2556])); 
mux_module mux_module_inst_1_2284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5111]),.i2(intermediate_reg_0[5110]),.o(intermediate_reg_1[2555]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5109]),.i2(intermediate_reg_0[5108]),.o(intermediate_reg_1[2554])); 
mux_module mux_module_inst_1_2286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5107]),.i2(intermediate_reg_0[5106]),.o(intermediate_reg_1[2553]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5105]),.i2(intermediate_reg_0[5104]),.o(intermediate_reg_1[2552])); 
mux_module mux_module_inst_1_2288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5103]),.i2(intermediate_reg_0[5102]),.o(intermediate_reg_1[2551]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5101]),.i2(intermediate_reg_0[5100]),.o(intermediate_reg_1[2550]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5099]),.i2(intermediate_reg_0[5098]),.o(intermediate_reg_1[2549])); 
mux_module mux_module_inst_1_2291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5097]),.i2(intermediate_reg_0[5096]),.o(intermediate_reg_1[2548]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5095]),.i2(intermediate_reg_0[5094]),.o(intermediate_reg_1[2547])); 
mux_module mux_module_inst_1_2293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5093]),.i2(intermediate_reg_0[5092]),.o(intermediate_reg_1[2546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5091]),.i2(intermediate_reg_0[5090]),.o(intermediate_reg_1[2545]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5089]),.i2(intermediate_reg_0[5088]),.o(intermediate_reg_1[2544])); 
mux_module mux_module_inst_1_2296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5087]),.i2(intermediate_reg_0[5086]),.o(intermediate_reg_1[2543]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5085]),.i2(intermediate_reg_0[5084]),.o(intermediate_reg_1[2542]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5083]),.i2(intermediate_reg_0[5082]),.o(intermediate_reg_1[2541])); 
mux_module mux_module_inst_1_2299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5081]),.i2(intermediate_reg_0[5080]),.o(intermediate_reg_1[2540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5079]),.i2(intermediate_reg_0[5078]),.o(intermediate_reg_1[2539]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5077]),.i2(intermediate_reg_0[5076]),.o(intermediate_reg_1[2538])); 
mux_module mux_module_inst_1_2302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5075]),.i2(intermediate_reg_0[5074]),.o(intermediate_reg_1[2537]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5073]),.i2(intermediate_reg_0[5072]),.o(intermediate_reg_1[2536])); 
fsm fsm_inst_1_2304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5071]),.i2(intermediate_reg_0[5070]),.o(intermediate_reg_1[2535])); 
fsm fsm_inst_1_2305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5069]),.i2(intermediate_reg_0[5068]),.o(intermediate_reg_1[2534])); 
mux_module mux_module_inst_1_2306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5067]),.i2(intermediate_reg_0[5066]),.o(intermediate_reg_1[2533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5065]),.i2(intermediate_reg_0[5064]),.o(intermediate_reg_1[2532]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5063]),.i2(intermediate_reg_0[5062]),.o(intermediate_reg_1[2531])); 
fsm fsm_inst_1_2309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5061]),.i2(intermediate_reg_0[5060]),.o(intermediate_reg_1[2530])); 
mux_module mux_module_inst_1_2310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5059]),.i2(intermediate_reg_0[5058]),.o(intermediate_reg_1[2529]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5057]),.i2(intermediate_reg_0[5056]),.o(intermediate_reg_1[2528])); 
fsm fsm_inst_1_2312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5055]),.i2(intermediate_reg_0[5054]),.o(intermediate_reg_1[2527])); 
mux_module mux_module_inst_1_2313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5053]),.i2(intermediate_reg_0[5052]),.o(intermediate_reg_1[2526]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5051]),.i2(intermediate_reg_0[5050]),.o(intermediate_reg_1[2525])); 
mux_module mux_module_inst_1_2315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5049]),.i2(intermediate_reg_0[5048]),.o(intermediate_reg_1[2524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5047]),.i2(intermediate_reg_0[5046]),.o(intermediate_reg_1[2523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5045]),.i2(intermediate_reg_0[5044]),.o(intermediate_reg_1[2522]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5043]),.i2(intermediate_reg_0[5042]),.o(intermediate_reg_1[2521])); 
mux_module mux_module_inst_1_2319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5041]),.i2(intermediate_reg_0[5040]),.o(intermediate_reg_1[2520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5039]),.i2(intermediate_reg_0[5038]),.o(intermediate_reg_1[2519]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5037]),.i2(intermediate_reg_0[5036]),.o(intermediate_reg_1[2518])); 
fsm fsm_inst_1_2322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5035]),.i2(intermediate_reg_0[5034]),.o(intermediate_reg_1[2517])); 
fsm fsm_inst_1_2323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5033]),.i2(intermediate_reg_0[5032]),.o(intermediate_reg_1[2516])); 
mux_module mux_module_inst_1_2324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5031]),.i2(intermediate_reg_0[5030]),.o(intermediate_reg_1[2515]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5029]),.i2(intermediate_reg_0[5028]),.o(intermediate_reg_1[2514])); 
fsm fsm_inst_1_2326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5027]),.i2(intermediate_reg_0[5026]),.o(intermediate_reg_1[2513])); 
mux_module mux_module_inst_1_2327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5025]),.i2(intermediate_reg_0[5024]),.o(intermediate_reg_1[2512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5023]),.i2(intermediate_reg_0[5022]),.o(intermediate_reg_1[2511]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5021]),.i2(intermediate_reg_0[5020]),.o(intermediate_reg_1[2510])); 
mux_module mux_module_inst_1_2330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5019]),.i2(intermediate_reg_0[5018]),.o(intermediate_reg_1[2509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5017]),.i2(intermediate_reg_0[5016]),.o(intermediate_reg_1[2508]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5015]),.i2(intermediate_reg_0[5014]),.o(intermediate_reg_1[2507]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5013]),.i2(intermediate_reg_0[5012]),.o(intermediate_reg_1[2506])); 
mux_module mux_module_inst_1_2334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5011]),.i2(intermediate_reg_0[5010]),.o(intermediate_reg_1[2505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5009]),.i2(intermediate_reg_0[5008]),.o(intermediate_reg_1[2504]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5007]),.i2(intermediate_reg_0[5006]),.o(intermediate_reg_1[2503]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5005]),.i2(intermediate_reg_0[5004]),.o(intermediate_reg_1[2502])); 
fsm fsm_inst_1_2338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5003]),.i2(intermediate_reg_0[5002]),.o(intermediate_reg_1[2501])); 
fsm fsm_inst_1_2339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5001]),.i2(intermediate_reg_0[5000]),.o(intermediate_reg_1[2500])); 
mux_module mux_module_inst_1_2340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4999]),.i2(intermediate_reg_0[4998]),.o(intermediate_reg_1[2499]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4997]),.i2(intermediate_reg_0[4996]),.o(intermediate_reg_1[2498])); 
fsm fsm_inst_1_2342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4995]),.i2(intermediate_reg_0[4994]),.o(intermediate_reg_1[2497])); 
fsm fsm_inst_1_2343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4993]),.i2(intermediate_reg_0[4992]),.o(intermediate_reg_1[2496])); 
mux_module mux_module_inst_1_2344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4991]),.i2(intermediate_reg_0[4990]),.o(intermediate_reg_1[2495]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4989]),.i2(intermediate_reg_0[4988]),.o(intermediate_reg_1[2494])); 
fsm fsm_inst_1_2346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4987]),.i2(intermediate_reg_0[4986]),.o(intermediate_reg_1[2493])); 
mux_module mux_module_inst_1_2347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4985]),.i2(intermediate_reg_0[4984]),.o(intermediate_reg_1[2492]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4983]),.i2(intermediate_reg_0[4982]),.o(intermediate_reg_1[2491])); 
mux_module mux_module_inst_1_2349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4981]),.i2(intermediate_reg_0[4980]),.o(intermediate_reg_1[2490]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4979]),.i2(intermediate_reg_0[4978]),.o(intermediate_reg_1[2489]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4977]),.i2(intermediate_reg_0[4976]),.o(intermediate_reg_1[2488]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4975]),.i2(intermediate_reg_0[4974]),.o(intermediate_reg_1[2487])); 
mux_module mux_module_inst_1_2353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4973]),.i2(intermediate_reg_0[4972]),.o(intermediate_reg_1[2486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4971]),.i2(intermediate_reg_0[4970]),.o(intermediate_reg_1[2485]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4969]),.i2(intermediate_reg_0[4968]),.o(intermediate_reg_1[2484])); 
fsm fsm_inst_1_2356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4967]),.i2(intermediate_reg_0[4966]),.o(intermediate_reg_1[2483])); 
mux_module mux_module_inst_1_2357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4965]),.i2(intermediate_reg_0[4964]),.o(intermediate_reg_1[2482]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4963]),.i2(intermediate_reg_0[4962]),.o(intermediate_reg_1[2481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4961]),.i2(intermediate_reg_0[4960]),.o(intermediate_reg_1[2480]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4959]),.i2(intermediate_reg_0[4958]),.o(intermediate_reg_1[2479]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4957]),.i2(intermediate_reg_0[4956]),.o(intermediate_reg_1[2478]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4955]),.i2(intermediate_reg_0[4954]),.o(intermediate_reg_1[2477])); 
mux_module mux_module_inst_1_2363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4953]),.i2(intermediate_reg_0[4952]),.o(intermediate_reg_1[2476]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4951]),.i2(intermediate_reg_0[4950]),.o(intermediate_reg_1[2475])); 
mux_module mux_module_inst_1_2365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4949]),.i2(intermediate_reg_0[4948]),.o(intermediate_reg_1[2474]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4947]),.i2(intermediate_reg_0[4946]),.o(intermediate_reg_1[2473])); 
fsm fsm_inst_1_2367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4945]),.i2(intermediate_reg_0[4944]),.o(intermediate_reg_1[2472])); 
mux_module mux_module_inst_1_2368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4943]),.i2(intermediate_reg_0[4942]),.o(intermediate_reg_1[2471]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4941]),.i2(intermediate_reg_0[4940]),.o(intermediate_reg_1[2470])); 
fsm fsm_inst_1_2370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4939]),.i2(intermediate_reg_0[4938]),.o(intermediate_reg_1[2469])); 
fsm fsm_inst_1_2371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4937]),.i2(intermediate_reg_0[4936]),.o(intermediate_reg_1[2468])); 
mux_module mux_module_inst_1_2372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4935]),.i2(intermediate_reg_0[4934]),.o(intermediate_reg_1[2467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4933]),.i2(intermediate_reg_0[4932]),.o(intermediate_reg_1[2466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4931]),.i2(intermediate_reg_0[4930]),.o(intermediate_reg_1[2465]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4929]),.i2(intermediate_reg_0[4928]),.o(intermediate_reg_1[2464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4927]),.i2(intermediate_reg_0[4926]),.o(intermediate_reg_1[2463]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4925]),.i2(intermediate_reg_0[4924]),.o(intermediate_reg_1[2462]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4923]),.i2(intermediate_reg_0[4922]),.o(intermediate_reg_1[2461])); 
mux_module mux_module_inst_1_2379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4921]),.i2(intermediate_reg_0[4920]),.o(intermediate_reg_1[2460]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4919]),.i2(intermediate_reg_0[4918]),.o(intermediate_reg_1[2459])); 
mux_module mux_module_inst_1_2381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4917]),.i2(intermediate_reg_0[4916]),.o(intermediate_reg_1[2458]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4915]),.i2(intermediate_reg_0[4914]),.o(intermediate_reg_1[2457])); 
fsm fsm_inst_1_2383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4913]),.i2(intermediate_reg_0[4912]),.o(intermediate_reg_1[2456])); 
fsm fsm_inst_1_2384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4911]),.i2(intermediate_reg_0[4910]),.o(intermediate_reg_1[2455])); 
mux_module mux_module_inst_1_2385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4909]),.i2(intermediate_reg_0[4908]),.o(intermediate_reg_1[2454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4907]),.i2(intermediate_reg_0[4906]),.o(intermediate_reg_1[2453]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4905]),.i2(intermediate_reg_0[4904]),.o(intermediate_reg_1[2452])); 
fsm fsm_inst_1_2388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4903]),.i2(intermediate_reg_0[4902]),.o(intermediate_reg_1[2451])); 
mux_module mux_module_inst_1_2389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4901]),.i2(intermediate_reg_0[4900]),.o(intermediate_reg_1[2450]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4899]),.i2(intermediate_reg_0[4898]),.o(intermediate_reg_1[2449])); 
mux_module mux_module_inst_1_2391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4897]),.i2(intermediate_reg_0[4896]),.o(intermediate_reg_1[2448]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4895]),.i2(intermediate_reg_0[4894]),.o(intermediate_reg_1[2447]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4893]),.i2(intermediate_reg_0[4892]),.o(intermediate_reg_1[2446]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4891]),.i2(intermediate_reg_0[4890]),.o(intermediate_reg_1[2445])); 
mux_module mux_module_inst_1_2395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4889]),.i2(intermediate_reg_0[4888]),.o(intermediate_reg_1[2444]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4887]),.i2(intermediate_reg_0[4886]),.o(intermediate_reg_1[2443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4885]),.i2(intermediate_reg_0[4884]),.o(intermediate_reg_1[2442]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4883]),.i2(intermediate_reg_0[4882]),.o(intermediate_reg_1[2441])); 
mux_module mux_module_inst_1_2399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4881]),.i2(intermediate_reg_0[4880]),.o(intermediate_reg_1[2440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4879]),.i2(intermediate_reg_0[4878]),.o(intermediate_reg_1[2439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4877]),.i2(intermediate_reg_0[4876]),.o(intermediate_reg_1[2438]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4875]),.i2(intermediate_reg_0[4874]),.o(intermediate_reg_1[2437])); 
mux_module mux_module_inst_1_2403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4873]),.i2(intermediate_reg_0[4872]),.o(intermediate_reg_1[2436]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4871]),.i2(intermediate_reg_0[4870]),.o(intermediate_reg_1[2435]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4869]),.i2(intermediate_reg_0[4868]),.o(intermediate_reg_1[2434]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4867]),.i2(intermediate_reg_0[4866]),.o(intermediate_reg_1[2433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4865]),.i2(intermediate_reg_0[4864]),.o(intermediate_reg_1[2432]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4863]),.i2(intermediate_reg_0[4862]),.o(intermediate_reg_1[2431])); 
mux_module mux_module_inst_1_2409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4861]),.i2(intermediate_reg_0[4860]),.o(intermediate_reg_1[2430]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4859]),.i2(intermediate_reg_0[4858]),.o(intermediate_reg_1[2429]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4857]),.i2(intermediate_reg_0[4856]),.o(intermediate_reg_1[2428])); 
mux_module mux_module_inst_1_2412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4855]),.i2(intermediate_reg_0[4854]),.o(intermediate_reg_1[2427]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4853]),.i2(intermediate_reg_0[4852]),.o(intermediate_reg_1[2426])); 
fsm fsm_inst_1_2414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4851]),.i2(intermediate_reg_0[4850]),.o(intermediate_reg_1[2425])); 
fsm fsm_inst_1_2415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4849]),.i2(intermediate_reg_0[4848]),.o(intermediate_reg_1[2424])); 
fsm fsm_inst_1_2416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4847]),.i2(intermediate_reg_0[4846]),.o(intermediate_reg_1[2423])); 
fsm fsm_inst_1_2417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4845]),.i2(intermediate_reg_0[4844]),.o(intermediate_reg_1[2422])); 
fsm fsm_inst_1_2418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4843]),.i2(intermediate_reg_0[4842]),.o(intermediate_reg_1[2421])); 
fsm fsm_inst_1_2419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4841]),.i2(intermediate_reg_0[4840]),.o(intermediate_reg_1[2420])); 
mux_module mux_module_inst_1_2420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4839]),.i2(intermediate_reg_0[4838]),.o(intermediate_reg_1[2419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4837]),.i2(intermediate_reg_0[4836]),.o(intermediate_reg_1[2418]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4835]),.i2(intermediate_reg_0[4834]),.o(intermediate_reg_1[2417]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4833]),.i2(intermediate_reg_0[4832]),.o(intermediate_reg_1[2416])); 
fsm fsm_inst_1_2424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4831]),.i2(intermediate_reg_0[4830]),.o(intermediate_reg_1[2415])); 
mux_module mux_module_inst_1_2425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4829]),.i2(intermediate_reg_0[4828]),.o(intermediate_reg_1[2414]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4827]),.i2(intermediate_reg_0[4826]),.o(intermediate_reg_1[2413]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4825]),.i2(intermediate_reg_0[4824]),.o(intermediate_reg_1[2412])); 
mux_module mux_module_inst_1_2428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4823]),.i2(intermediate_reg_0[4822]),.o(intermediate_reg_1[2411]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4821]),.i2(intermediate_reg_0[4820]),.o(intermediate_reg_1[2410]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4819]),.i2(intermediate_reg_0[4818]),.o(intermediate_reg_1[2409]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4817]),.i2(intermediate_reg_0[4816]),.o(intermediate_reg_1[2408]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4815]),.i2(intermediate_reg_0[4814]),.o(intermediate_reg_1[2407])); 
mux_module mux_module_inst_1_2433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4813]),.i2(intermediate_reg_0[4812]),.o(intermediate_reg_1[2406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4811]),.i2(intermediate_reg_0[4810]),.o(intermediate_reg_1[2405]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4809]),.i2(intermediate_reg_0[4808]),.o(intermediate_reg_1[2404])); 
fsm fsm_inst_1_2436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4807]),.i2(intermediate_reg_0[4806]),.o(intermediate_reg_1[2403])); 
fsm fsm_inst_1_2437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4805]),.i2(intermediate_reg_0[4804]),.o(intermediate_reg_1[2402])); 
mux_module mux_module_inst_1_2438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4803]),.i2(intermediate_reg_0[4802]),.o(intermediate_reg_1[2401]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4801]),.i2(intermediate_reg_0[4800]),.o(intermediate_reg_1[2400])); 
fsm fsm_inst_1_2440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4799]),.i2(intermediate_reg_0[4798]),.o(intermediate_reg_1[2399])); 
mux_module mux_module_inst_1_2441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4797]),.i2(intermediate_reg_0[4796]),.o(intermediate_reg_1[2398]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4795]),.i2(intermediate_reg_0[4794]),.o(intermediate_reg_1[2397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4793]),.i2(intermediate_reg_0[4792]),.o(intermediate_reg_1[2396]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4791]),.i2(intermediate_reg_0[4790]),.o(intermediate_reg_1[2395])); 
mux_module mux_module_inst_1_2445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4789]),.i2(intermediate_reg_0[4788]),.o(intermediate_reg_1[2394]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4787]),.i2(intermediate_reg_0[4786]),.o(intermediate_reg_1[2393])); 
mux_module mux_module_inst_1_2447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4785]),.i2(intermediate_reg_0[4784]),.o(intermediate_reg_1[2392]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4783]),.i2(intermediate_reg_0[4782]),.o(intermediate_reg_1[2391])); 
mux_module mux_module_inst_1_2449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4781]),.i2(intermediate_reg_0[4780]),.o(intermediate_reg_1[2390]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4779]),.i2(intermediate_reg_0[4778]),.o(intermediate_reg_1[2389])); 
mux_module mux_module_inst_1_2451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4777]),.i2(intermediate_reg_0[4776]),.o(intermediate_reg_1[2388]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4775]),.i2(intermediate_reg_0[4774]),.o(intermediate_reg_1[2387])); 
mux_module mux_module_inst_1_2453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4773]),.i2(intermediate_reg_0[4772]),.o(intermediate_reg_1[2386]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4771]),.i2(intermediate_reg_0[4770]),.o(intermediate_reg_1[2385]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4769]),.i2(intermediate_reg_0[4768]),.o(intermediate_reg_1[2384])); 
mux_module mux_module_inst_1_2456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4767]),.i2(intermediate_reg_0[4766]),.o(intermediate_reg_1[2383]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4765]),.i2(intermediate_reg_0[4764]),.o(intermediate_reg_1[2382])); 
fsm fsm_inst_1_2458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4763]),.i2(intermediate_reg_0[4762]),.o(intermediate_reg_1[2381])); 
fsm fsm_inst_1_2459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4761]),.i2(intermediate_reg_0[4760]),.o(intermediate_reg_1[2380])); 
fsm fsm_inst_1_2460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4759]),.i2(intermediate_reg_0[4758]),.o(intermediate_reg_1[2379])); 
fsm fsm_inst_1_2461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4757]),.i2(intermediate_reg_0[4756]),.o(intermediate_reg_1[2378])); 
fsm fsm_inst_1_2462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4755]),.i2(intermediate_reg_0[4754]),.o(intermediate_reg_1[2377])); 
mux_module mux_module_inst_1_2463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4753]),.i2(intermediate_reg_0[4752]),.o(intermediate_reg_1[2376]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4751]),.i2(intermediate_reg_0[4750]),.o(intermediate_reg_1[2375]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4749]),.i2(intermediate_reg_0[4748]),.o(intermediate_reg_1[2374])); 
fsm fsm_inst_1_2466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4747]),.i2(intermediate_reg_0[4746]),.o(intermediate_reg_1[2373])); 
mux_module mux_module_inst_1_2467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4745]),.i2(intermediate_reg_0[4744]),.o(intermediate_reg_1[2372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4743]),.i2(intermediate_reg_0[4742]),.o(intermediate_reg_1[2371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4741]),.i2(intermediate_reg_0[4740]),.o(intermediate_reg_1[2370]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4739]),.i2(intermediate_reg_0[4738]),.o(intermediate_reg_1[2369])); 
mux_module mux_module_inst_1_2471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4737]),.i2(intermediate_reg_0[4736]),.o(intermediate_reg_1[2368]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4735]),.i2(intermediate_reg_0[4734]),.o(intermediate_reg_1[2367])); 
fsm fsm_inst_1_2473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4733]),.i2(intermediate_reg_0[4732]),.o(intermediate_reg_1[2366])); 
fsm fsm_inst_1_2474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4731]),.i2(intermediate_reg_0[4730]),.o(intermediate_reg_1[2365])); 
mux_module mux_module_inst_1_2475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4729]),.i2(intermediate_reg_0[4728]),.o(intermediate_reg_1[2364]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4727]),.i2(intermediate_reg_0[4726]),.o(intermediate_reg_1[2363]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4725]),.i2(intermediate_reg_0[4724]),.o(intermediate_reg_1[2362])); 
fsm fsm_inst_1_2478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4723]),.i2(intermediate_reg_0[4722]),.o(intermediate_reg_1[2361])); 
fsm fsm_inst_1_2479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4721]),.i2(intermediate_reg_0[4720]),.o(intermediate_reg_1[2360])); 
mux_module mux_module_inst_1_2480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4719]),.i2(intermediate_reg_0[4718]),.o(intermediate_reg_1[2359]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4717]),.i2(intermediate_reg_0[4716]),.o(intermediate_reg_1[2358])); 
fsm fsm_inst_1_2482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4715]),.i2(intermediate_reg_0[4714]),.o(intermediate_reg_1[2357])); 
mux_module mux_module_inst_1_2483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4713]),.i2(intermediate_reg_0[4712]),.o(intermediate_reg_1[2356]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4711]),.i2(intermediate_reg_0[4710]),.o(intermediate_reg_1[2355]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4709]),.i2(intermediate_reg_0[4708]),.o(intermediate_reg_1[2354])); 
fsm fsm_inst_1_2486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4707]),.i2(intermediate_reg_0[4706]),.o(intermediate_reg_1[2353])); 
mux_module mux_module_inst_1_2487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4705]),.i2(intermediate_reg_0[4704]),.o(intermediate_reg_1[2352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4703]),.i2(intermediate_reg_0[4702]),.o(intermediate_reg_1[2351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4701]),.i2(intermediate_reg_0[4700]),.o(intermediate_reg_1[2350]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4699]),.i2(intermediate_reg_0[4698]),.o(intermediate_reg_1[2349]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4697]),.i2(intermediate_reg_0[4696]),.o(intermediate_reg_1[2348])); 
fsm fsm_inst_1_2492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4695]),.i2(intermediate_reg_0[4694]),.o(intermediate_reg_1[2347])); 
fsm fsm_inst_1_2493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4693]),.i2(intermediate_reg_0[4692]),.o(intermediate_reg_1[2346])); 
fsm fsm_inst_1_2494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4691]),.i2(intermediate_reg_0[4690]),.o(intermediate_reg_1[2345])); 
mux_module mux_module_inst_1_2495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4689]),.i2(intermediate_reg_0[4688]),.o(intermediate_reg_1[2344]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4687]),.i2(intermediate_reg_0[4686]),.o(intermediate_reg_1[2343]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4685]),.i2(intermediate_reg_0[4684]),.o(intermediate_reg_1[2342]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4683]),.i2(intermediate_reg_0[4682]),.o(intermediate_reg_1[2341])); 
mux_module mux_module_inst_1_2499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4681]),.i2(intermediate_reg_0[4680]),.o(intermediate_reg_1[2340]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4679]),.i2(intermediate_reg_0[4678]),.o(intermediate_reg_1[2339])); 
mux_module mux_module_inst_1_2501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4677]),.i2(intermediate_reg_0[4676]),.o(intermediate_reg_1[2338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4675]),.i2(intermediate_reg_0[4674]),.o(intermediate_reg_1[2337]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4673]),.i2(intermediate_reg_0[4672]),.o(intermediate_reg_1[2336])); 
fsm fsm_inst_1_2504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4671]),.i2(intermediate_reg_0[4670]),.o(intermediate_reg_1[2335])); 
fsm fsm_inst_1_2505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4669]),.i2(intermediate_reg_0[4668]),.o(intermediate_reg_1[2334])); 
mux_module mux_module_inst_1_2506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4667]),.i2(intermediate_reg_0[4666]),.o(intermediate_reg_1[2333]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4665]),.i2(intermediate_reg_0[4664]),.o(intermediate_reg_1[2332]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4663]),.i2(intermediate_reg_0[4662]),.o(intermediate_reg_1[2331])); 
mux_module mux_module_inst_1_2509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4661]),.i2(intermediate_reg_0[4660]),.o(intermediate_reg_1[2330]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4659]),.i2(intermediate_reg_0[4658]),.o(intermediate_reg_1[2329])); 
mux_module mux_module_inst_1_2511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4657]),.i2(intermediate_reg_0[4656]),.o(intermediate_reg_1[2328]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4655]),.i2(intermediate_reg_0[4654]),.o(intermediate_reg_1[2327])); 
fsm fsm_inst_1_2513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4653]),.i2(intermediate_reg_0[4652]),.o(intermediate_reg_1[2326])); 
fsm fsm_inst_1_2514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4651]),.i2(intermediate_reg_0[4650]),.o(intermediate_reg_1[2325])); 
mux_module mux_module_inst_1_2515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4649]),.i2(intermediate_reg_0[4648]),.o(intermediate_reg_1[2324]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4647]),.i2(intermediate_reg_0[4646]),.o(intermediate_reg_1[2323])); 
mux_module mux_module_inst_1_2517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4645]),.i2(intermediate_reg_0[4644]),.o(intermediate_reg_1[2322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4643]),.i2(intermediate_reg_0[4642]),.o(intermediate_reg_1[2321]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4641]),.i2(intermediate_reg_0[4640]),.o(intermediate_reg_1[2320])); 
mux_module mux_module_inst_1_2520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4639]),.i2(intermediate_reg_0[4638]),.o(intermediate_reg_1[2319]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4637]),.i2(intermediate_reg_0[4636]),.o(intermediate_reg_1[2318])); 
fsm fsm_inst_1_2522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4635]),.i2(intermediate_reg_0[4634]),.o(intermediate_reg_1[2317])); 
mux_module mux_module_inst_1_2523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4633]),.i2(intermediate_reg_0[4632]),.o(intermediate_reg_1[2316]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4631]),.i2(intermediate_reg_0[4630]),.o(intermediate_reg_1[2315])); 
mux_module mux_module_inst_1_2525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4629]),.i2(intermediate_reg_0[4628]),.o(intermediate_reg_1[2314]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4627]),.i2(intermediate_reg_0[4626]),.o(intermediate_reg_1[2313])); 
mux_module mux_module_inst_1_2527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4625]),.i2(intermediate_reg_0[4624]),.o(intermediate_reg_1[2312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4623]),.i2(intermediate_reg_0[4622]),.o(intermediate_reg_1[2311]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4621]),.i2(intermediate_reg_0[4620]),.o(intermediate_reg_1[2310])); 
fsm fsm_inst_1_2530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4619]),.i2(intermediate_reg_0[4618]),.o(intermediate_reg_1[2309])); 
fsm fsm_inst_1_2531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4617]),.i2(intermediate_reg_0[4616]),.o(intermediate_reg_1[2308])); 
fsm fsm_inst_1_2532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4615]),.i2(intermediate_reg_0[4614]),.o(intermediate_reg_1[2307])); 
fsm fsm_inst_1_2533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4613]),.i2(intermediate_reg_0[4612]),.o(intermediate_reg_1[2306])); 
mux_module mux_module_inst_1_2534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4611]),.i2(intermediate_reg_0[4610]),.o(intermediate_reg_1[2305]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4609]),.i2(intermediate_reg_0[4608]),.o(intermediate_reg_1[2304])); 
fsm fsm_inst_1_2536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4607]),.i2(intermediate_reg_0[4606]),.o(intermediate_reg_1[2303])); 
fsm fsm_inst_1_2537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4605]),.i2(intermediate_reg_0[4604]),.o(intermediate_reg_1[2302])); 
mux_module mux_module_inst_1_2538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4603]),.i2(intermediate_reg_0[4602]),.o(intermediate_reg_1[2301]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4601]),.i2(intermediate_reg_0[4600]),.o(intermediate_reg_1[2300])); 
fsm fsm_inst_1_2540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4599]),.i2(intermediate_reg_0[4598]),.o(intermediate_reg_1[2299])); 
mux_module mux_module_inst_1_2541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4597]),.i2(intermediate_reg_0[4596]),.o(intermediate_reg_1[2298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4595]),.i2(intermediate_reg_0[4594]),.o(intermediate_reg_1[2297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4593]),.i2(intermediate_reg_0[4592]),.o(intermediate_reg_1[2296]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4591]),.i2(intermediate_reg_0[4590]),.o(intermediate_reg_1[2295])); 
fsm fsm_inst_1_2545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4589]),.i2(intermediate_reg_0[4588]),.o(intermediate_reg_1[2294])); 
mux_module mux_module_inst_1_2546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4587]),.i2(intermediate_reg_0[4586]),.o(intermediate_reg_1[2293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4585]),.i2(intermediate_reg_0[4584]),.o(intermediate_reg_1[2292]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4583]),.i2(intermediate_reg_0[4582]),.o(intermediate_reg_1[2291])); 
fsm fsm_inst_1_2549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4581]),.i2(intermediate_reg_0[4580]),.o(intermediate_reg_1[2290])); 
mux_module mux_module_inst_1_2550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4579]),.i2(intermediate_reg_0[4578]),.o(intermediate_reg_1[2289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4577]),.i2(intermediate_reg_0[4576]),.o(intermediate_reg_1[2288]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4575]),.i2(intermediate_reg_0[4574]),.o(intermediate_reg_1[2287])); 
fsm fsm_inst_1_2553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4573]),.i2(intermediate_reg_0[4572]),.o(intermediate_reg_1[2286])); 
fsm fsm_inst_1_2554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4571]),.i2(intermediate_reg_0[4570]),.o(intermediate_reg_1[2285])); 
mux_module mux_module_inst_1_2555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4569]),.i2(intermediate_reg_0[4568]),.o(intermediate_reg_1[2284]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4567]),.i2(intermediate_reg_0[4566]),.o(intermediate_reg_1[2283])); 
mux_module mux_module_inst_1_2557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4565]),.i2(intermediate_reg_0[4564]),.o(intermediate_reg_1[2282]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4563]),.i2(intermediate_reg_0[4562]),.o(intermediate_reg_1[2281])); 
mux_module mux_module_inst_1_2559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4561]),.i2(intermediate_reg_0[4560]),.o(intermediate_reg_1[2280]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4559]),.i2(intermediate_reg_0[4558]),.o(intermediate_reg_1[2279]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4557]),.i2(intermediate_reg_0[4556]),.o(intermediate_reg_1[2278])); 
mux_module mux_module_inst_1_2562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4555]),.i2(intermediate_reg_0[4554]),.o(intermediate_reg_1[2277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4553]),.i2(intermediate_reg_0[4552]),.o(intermediate_reg_1[2276]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4551]),.i2(intermediate_reg_0[4550]),.o(intermediate_reg_1[2275])); 
mux_module mux_module_inst_1_2565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4549]),.i2(intermediate_reg_0[4548]),.o(intermediate_reg_1[2274]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4547]),.i2(intermediate_reg_0[4546]),.o(intermediate_reg_1[2273]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4545]),.i2(intermediate_reg_0[4544]),.o(intermediate_reg_1[2272]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4543]),.i2(intermediate_reg_0[4542]),.o(intermediate_reg_1[2271])); 
fsm fsm_inst_1_2569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4541]),.i2(intermediate_reg_0[4540]),.o(intermediate_reg_1[2270])); 
mux_module mux_module_inst_1_2570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4539]),.i2(intermediate_reg_0[4538]),.o(intermediate_reg_1[2269]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4537]),.i2(intermediate_reg_0[4536]),.o(intermediate_reg_1[2268])); 
fsm fsm_inst_1_2572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4535]),.i2(intermediate_reg_0[4534]),.o(intermediate_reg_1[2267])); 
mux_module mux_module_inst_1_2573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4533]),.i2(intermediate_reg_0[4532]),.o(intermediate_reg_1[2266]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4531]),.i2(intermediate_reg_0[4530]),.o(intermediate_reg_1[2265])); 
mux_module mux_module_inst_1_2575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4529]),.i2(intermediate_reg_0[4528]),.o(intermediate_reg_1[2264]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4527]),.i2(intermediate_reg_0[4526]),.o(intermediate_reg_1[2263])); 
mux_module mux_module_inst_1_2577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4525]),.i2(intermediate_reg_0[4524]),.o(intermediate_reg_1[2262]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4523]),.i2(intermediate_reg_0[4522]),.o(intermediate_reg_1[2261])); 
mux_module mux_module_inst_1_2579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4521]),.i2(intermediate_reg_0[4520]),.o(intermediate_reg_1[2260]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4519]),.i2(intermediate_reg_0[4518]),.o(intermediate_reg_1[2259])); 
fsm fsm_inst_1_2581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4517]),.i2(intermediate_reg_0[4516]),.o(intermediate_reg_1[2258])); 
mux_module mux_module_inst_1_2582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4515]),.i2(intermediate_reg_0[4514]),.o(intermediate_reg_1[2257]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4513]),.i2(intermediate_reg_0[4512]),.o(intermediate_reg_1[2256])); 
mux_module mux_module_inst_1_2584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4511]),.i2(intermediate_reg_0[4510]),.o(intermediate_reg_1[2255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4509]),.i2(intermediate_reg_0[4508]),.o(intermediate_reg_1[2254]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4507]),.i2(intermediate_reg_0[4506]),.o(intermediate_reg_1[2253])); 
fsm fsm_inst_1_2587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4505]),.i2(intermediate_reg_0[4504]),.o(intermediate_reg_1[2252])); 
fsm fsm_inst_1_2588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4503]),.i2(intermediate_reg_0[4502]),.o(intermediate_reg_1[2251])); 
mux_module mux_module_inst_1_2589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4501]),.i2(intermediate_reg_0[4500]),.o(intermediate_reg_1[2250]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4499]),.i2(intermediate_reg_0[4498]),.o(intermediate_reg_1[2249])); 
mux_module mux_module_inst_1_2591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4497]),.i2(intermediate_reg_0[4496]),.o(intermediate_reg_1[2248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4495]),.i2(intermediate_reg_0[4494]),.o(intermediate_reg_1[2247]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4493]),.i2(intermediate_reg_0[4492]),.o(intermediate_reg_1[2246])); 
fsm fsm_inst_1_2594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4491]),.i2(intermediate_reg_0[4490]),.o(intermediate_reg_1[2245])); 
mux_module mux_module_inst_1_2595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4489]),.i2(intermediate_reg_0[4488]),.o(intermediate_reg_1[2244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4487]),.i2(intermediate_reg_0[4486]),.o(intermediate_reg_1[2243]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4485]),.i2(intermediate_reg_0[4484]),.o(intermediate_reg_1[2242]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4483]),.i2(intermediate_reg_0[4482]),.o(intermediate_reg_1[2241])); 
mux_module mux_module_inst_1_2599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4481]),.i2(intermediate_reg_0[4480]),.o(intermediate_reg_1[2240]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4479]),.i2(intermediate_reg_0[4478]),.o(intermediate_reg_1[2239])); 
fsm fsm_inst_1_2601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4477]),.i2(intermediate_reg_0[4476]),.o(intermediate_reg_1[2238])); 
mux_module mux_module_inst_1_2602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4475]),.i2(intermediate_reg_0[4474]),.o(intermediate_reg_1[2237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4473]),.i2(intermediate_reg_0[4472]),.o(intermediate_reg_1[2236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4471]),.i2(intermediate_reg_0[4470]),.o(intermediate_reg_1[2235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4469]),.i2(intermediate_reg_0[4468]),.o(intermediate_reg_1[2234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4467]),.i2(intermediate_reg_0[4466]),.o(intermediate_reg_1[2233]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4465]),.i2(intermediate_reg_0[4464]),.o(intermediate_reg_1[2232]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4463]),.i2(intermediate_reg_0[4462]),.o(intermediate_reg_1[2231])); 
fsm fsm_inst_1_2609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4461]),.i2(intermediate_reg_0[4460]),.o(intermediate_reg_1[2230])); 
mux_module mux_module_inst_1_2610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4459]),.i2(intermediate_reg_0[4458]),.o(intermediate_reg_1[2229]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4457]),.i2(intermediate_reg_0[4456]),.o(intermediate_reg_1[2228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4455]),.i2(intermediate_reg_0[4454]),.o(intermediate_reg_1[2227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4453]),.i2(intermediate_reg_0[4452]),.o(intermediate_reg_1[2226]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4451]),.i2(intermediate_reg_0[4450]),.o(intermediate_reg_1[2225])); 
fsm fsm_inst_1_2615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4449]),.i2(intermediate_reg_0[4448]),.o(intermediate_reg_1[2224])); 
fsm fsm_inst_1_2616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4447]),.i2(intermediate_reg_0[4446]),.o(intermediate_reg_1[2223])); 
fsm fsm_inst_1_2617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4445]),.i2(intermediate_reg_0[4444]),.o(intermediate_reg_1[2222])); 
mux_module mux_module_inst_1_2618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4443]),.i2(intermediate_reg_0[4442]),.o(intermediate_reg_1[2221]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4441]),.i2(intermediate_reg_0[4440]),.o(intermediate_reg_1[2220])); 
mux_module mux_module_inst_1_2620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4439]),.i2(intermediate_reg_0[4438]),.o(intermediate_reg_1[2219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4437]),.i2(intermediate_reg_0[4436]),.o(intermediate_reg_1[2218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4435]),.i2(intermediate_reg_0[4434]),.o(intermediate_reg_1[2217]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4433]),.i2(intermediate_reg_0[4432]),.o(intermediate_reg_1[2216])); 
fsm fsm_inst_1_2624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4431]),.i2(intermediate_reg_0[4430]),.o(intermediate_reg_1[2215])); 
mux_module mux_module_inst_1_2625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4429]),.i2(intermediate_reg_0[4428]),.o(intermediate_reg_1[2214]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4427]),.i2(intermediate_reg_0[4426]),.o(intermediate_reg_1[2213])); 
fsm fsm_inst_1_2627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4425]),.i2(intermediate_reg_0[4424]),.o(intermediate_reg_1[2212])); 
mux_module mux_module_inst_1_2628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4423]),.i2(intermediate_reg_0[4422]),.o(intermediate_reg_1[2211]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4421]),.i2(intermediate_reg_0[4420]),.o(intermediate_reg_1[2210])); 
fsm fsm_inst_1_2630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4419]),.i2(intermediate_reg_0[4418]),.o(intermediate_reg_1[2209])); 
fsm fsm_inst_1_2631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4417]),.i2(intermediate_reg_0[4416]),.o(intermediate_reg_1[2208])); 
fsm fsm_inst_1_2632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4415]),.i2(intermediate_reg_0[4414]),.o(intermediate_reg_1[2207])); 
fsm fsm_inst_1_2633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4413]),.i2(intermediate_reg_0[4412]),.o(intermediate_reg_1[2206])); 
mux_module mux_module_inst_1_2634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4411]),.i2(intermediate_reg_0[4410]),.o(intermediate_reg_1[2205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4409]),.i2(intermediate_reg_0[4408]),.o(intermediate_reg_1[2204]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4407]),.i2(intermediate_reg_0[4406]),.o(intermediate_reg_1[2203])); 
mux_module mux_module_inst_1_2637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4405]),.i2(intermediate_reg_0[4404]),.o(intermediate_reg_1[2202]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4403]),.i2(intermediate_reg_0[4402]),.o(intermediate_reg_1[2201]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4401]),.i2(intermediate_reg_0[4400]),.o(intermediate_reg_1[2200])); 
fsm fsm_inst_1_2640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4399]),.i2(intermediate_reg_0[4398]),.o(intermediate_reg_1[2199])); 
mux_module mux_module_inst_1_2641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4397]),.i2(intermediate_reg_0[4396]),.o(intermediate_reg_1[2198]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4395]),.i2(intermediate_reg_0[4394]),.o(intermediate_reg_1[2197])); 
fsm fsm_inst_1_2643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4393]),.i2(intermediate_reg_0[4392]),.o(intermediate_reg_1[2196])); 
fsm fsm_inst_1_2644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4391]),.i2(intermediate_reg_0[4390]),.o(intermediate_reg_1[2195])); 
mux_module mux_module_inst_1_2645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4389]),.i2(intermediate_reg_0[4388]),.o(intermediate_reg_1[2194]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4387]),.i2(intermediate_reg_0[4386]),.o(intermediate_reg_1[2193])); 
fsm fsm_inst_1_2647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4385]),.i2(intermediate_reg_0[4384]),.o(intermediate_reg_1[2192])); 
fsm fsm_inst_1_2648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4383]),.i2(intermediate_reg_0[4382]),.o(intermediate_reg_1[2191])); 
mux_module mux_module_inst_1_2649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4381]),.i2(intermediate_reg_0[4380]),.o(intermediate_reg_1[2190]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4379]),.i2(intermediate_reg_0[4378]),.o(intermediate_reg_1[2189])); 
mux_module mux_module_inst_1_2651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4377]),.i2(intermediate_reg_0[4376]),.o(intermediate_reg_1[2188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4375]),.i2(intermediate_reg_0[4374]),.o(intermediate_reg_1[2187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4373]),.i2(intermediate_reg_0[4372]),.o(intermediate_reg_1[2186]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4371]),.i2(intermediate_reg_0[4370]),.o(intermediate_reg_1[2185])); 
fsm fsm_inst_1_2655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4369]),.i2(intermediate_reg_0[4368]),.o(intermediate_reg_1[2184])); 
mux_module mux_module_inst_1_2656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4367]),.i2(intermediate_reg_0[4366]),.o(intermediate_reg_1[2183]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4365]),.i2(intermediate_reg_0[4364]),.o(intermediate_reg_1[2182])); 
mux_module mux_module_inst_1_2658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4363]),.i2(intermediate_reg_0[4362]),.o(intermediate_reg_1[2181]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4361]),.i2(intermediate_reg_0[4360]),.o(intermediate_reg_1[2180])); 
mux_module mux_module_inst_1_2660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4359]),.i2(intermediate_reg_0[4358]),.o(intermediate_reg_1[2179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4357]),.i2(intermediate_reg_0[4356]),.o(intermediate_reg_1[2178]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4355]),.i2(intermediate_reg_0[4354]),.o(intermediate_reg_1[2177])); 
fsm fsm_inst_1_2663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4353]),.i2(intermediate_reg_0[4352]),.o(intermediate_reg_1[2176])); 
fsm fsm_inst_1_2664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4351]),.i2(intermediate_reg_0[4350]),.o(intermediate_reg_1[2175])); 
mux_module mux_module_inst_1_2665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4349]),.i2(intermediate_reg_0[4348]),.o(intermediate_reg_1[2174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4347]),.i2(intermediate_reg_0[4346]),.o(intermediate_reg_1[2173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4345]),.i2(intermediate_reg_0[4344]),.o(intermediate_reg_1[2172]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4343]),.i2(intermediate_reg_0[4342]),.o(intermediate_reg_1[2171])); 
mux_module mux_module_inst_1_2669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4341]),.i2(intermediate_reg_0[4340]),.o(intermediate_reg_1[2170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4339]),.i2(intermediate_reg_0[4338]),.o(intermediate_reg_1[2169]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4337]),.i2(intermediate_reg_0[4336]),.o(intermediate_reg_1[2168])); 
mux_module mux_module_inst_1_2672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4335]),.i2(intermediate_reg_0[4334]),.o(intermediate_reg_1[2167]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4333]),.i2(intermediate_reg_0[4332]),.o(intermediate_reg_1[2166])); 
mux_module mux_module_inst_1_2674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4331]),.i2(intermediate_reg_0[4330]),.o(intermediate_reg_1[2165]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4329]),.i2(intermediate_reg_0[4328]),.o(intermediate_reg_1[2164])); 
mux_module mux_module_inst_1_2676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4327]),.i2(intermediate_reg_0[4326]),.o(intermediate_reg_1[2163]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4325]),.i2(intermediate_reg_0[4324]),.o(intermediate_reg_1[2162])); 
fsm fsm_inst_1_2678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4323]),.i2(intermediate_reg_0[4322]),.o(intermediate_reg_1[2161])); 
fsm fsm_inst_1_2679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4321]),.i2(intermediate_reg_0[4320]),.o(intermediate_reg_1[2160])); 
mux_module mux_module_inst_1_2680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4319]),.i2(intermediate_reg_0[4318]),.o(intermediate_reg_1[2159]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4317]),.i2(intermediate_reg_0[4316]),.o(intermediate_reg_1[2158])); 
mux_module mux_module_inst_1_2682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4315]),.i2(intermediate_reg_0[4314]),.o(intermediate_reg_1[2157]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4313]),.i2(intermediate_reg_0[4312]),.o(intermediate_reg_1[2156])); 
fsm fsm_inst_1_2684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4311]),.i2(intermediate_reg_0[4310]),.o(intermediate_reg_1[2155])); 
mux_module mux_module_inst_1_2685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4309]),.i2(intermediate_reg_0[4308]),.o(intermediate_reg_1[2154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4307]),.i2(intermediate_reg_0[4306]),.o(intermediate_reg_1[2153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4305]),.i2(intermediate_reg_0[4304]),.o(intermediate_reg_1[2152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4303]),.i2(intermediate_reg_0[4302]),.o(intermediate_reg_1[2151]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4301]),.i2(intermediate_reg_0[4300]),.o(intermediate_reg_1[2150])); 
mux_module mux_module_inst_1_2690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4299]),.i2(intermediate_reg_0[4298]),.o(intermediate_reg_1[2149]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4297]),.i2(intermediate_reg_0[4296]),.o(intermediate_reg_1[2148])); 
fsm fsm_inst_1_2692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4295]),.i2(intermediate_reg_0[4294]),.o(intermediate_reg_1[2147])); 
mux_module mux_module_inst_1_2693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4293]),.i2(intermediate_reg_0[4292]),.o(intermediate_reg_1[2146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4291]),.i2(intermediate_reg_0[4290]),.o(intermediate_reg_1[2145]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4289]),.i2(intermediate_reg_0[4288]),.o(intermediate_reg_1[2144])); 
fsm fsm_inst_1_2696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4287]),.i2(intermediate_reg_0[4286]),.o(intermediate_reg_1[2143])); 
mux_module mux_module_inst_1_2697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4285]),.i2(intermediate_reg_0[4284]),.o(intermediate_reg_1[2142]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4283]),.i2(intermediate_reg_0[4282]),.o(intermediate_reg_1[2141]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4281]),.i2(intermediate_reg_0[4280]),.o(intermediate_reg_1[2140])); 
mux_module mux_module_inst_1_2700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4279]),.i2(intermediate_reg_0[4278]),.o(intermediate_reg_1[2139]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4277]),.i2(intermediate_reg_0[4276]),.o(intermediate_reg_1[2138])); 
fsm fsm_inst_1_2702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4275]),.i2(intermediate_reg_0[4274]),.o(intermediate_reg_1[2137])); 
fsm fsm_inst_1_2703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4273]),.i2(intermediate_reg_0[4272]),.o(intermediate_reg_1[2136])); 
fsm fsm_inst_1_2704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4271]),.i2(intermediate_reg_0[4270]),.o(intermediate_reg_1[2135])); 
mux_module mux_module_inst_1_2705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4269]),.i2(intermediate_reg_0[4268]),.o(intermediate_reg_1[2134]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4267]),.i2(intermediate_reg_0[4266]),.o(intermediate_reg_1[2133]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4265]),.i2(intermediate_reg_0[4264]),.o(intermediate_reg_1[2132])); 
fsm fsm_inst_1_2708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4263]),.i2(intermediate_reg_0[4262]),.o(intermediate_reg_1[2131])); 
fsm fsm_inst_1_2709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4261]),.i2(intermediate_reg_0[4260]),.o(intermediate_reg_1[2130])); 
fsm fsm_inst_1_2710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4259]),.i2(intermediate_reg_0[4258]),.o(intermediate_reg_1[2129])); 
fsm fsm_inst_1_2711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4257]),.i2(intermediate_reg_0[4256]),.o(intermediate_reg_1[2128])); 
mux_module mux_module_inst_1_2712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4255]),.i2(intermediate_reg_0[4254]),.o(intermediate_reg_1[2127]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4253]),.i2(intermediate_reg_0[4252]),.o(intermediate_reg_1[2126])); 
fsm fsm_inst_1_2714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4251]),.i2(intermediate_reg_0[4250]),.o(intermediate_reg_1[2125])); 
fsm fsm_inst_1_2715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4249]),.i2(intermediate_reg_0[4248]),.o(intermediate_reg_1[2124])); 
fsm fsm_inst_1_2716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4247]),.i2(intermediate_reg_0[4246]),.o(intermediate_reg_1[2123])); 
fsm fsm_inst_1_2717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4245]),.i2(intermediate_reg_0[4244]),.o(intermediate_reg_1[2122])); 
fsm fsm_inst_1_2718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4243]),.i2(intermediate_reg_0[4242]),.o(intermediate_reg_1[2121])); 
mux_module mux_module_inst_1_2719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4241]),.i2(intermediate_reg_0[4240]),.o(intermediate_reg_1[2120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4239]),.i2(intermediate_reg_0[4238]),.o(intermediate_reg_1[2119]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4237]),.i2(intermediate_reg_0[4236]),.o(intermediate_reg_1[2118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4235]),.i2(intermediate_reg_0[4234]),.o(intermediate_reg_1[2117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4233]),.i2(intermediate_reg_0[4232]),.o(intermediate_reg_1[2116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4231]),.i2(intermediate_reg_0[4230]),.o(intermediate_reg_1[2115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4229]),.i2(intermediate_reg_0[4228]),.o(intermediate_reg_1[2114])); 
mux_module mux_module_inst_1_2726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4227]),.i2(intermediate_reg_0[4226]),.o(intermediate_reg_1[2113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4225]),.i2(intermediate_reg_0[4224]),.o(intermediate_reg_1[2112]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4223]),.i2(intermediate_reg_0[4222]),.o(intermediate_reg_1[2111])); 
fsm fsm_inst_1_2729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4221]),.i2(intermediate_reg_0[4220]),.o(intermediate_reg_1[2110])); 
mux_module mux_module_inst_1_2730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4219]),.i2(intermediate_reg_0[4218]),.o(intermediate_reg_1[2109]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4217]),.i2(intermediate_reg_0[4216]),.o(intermediate_reg_1[2108])); 
fsm fsm_inst_1_2732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4215]),.i2(intermediate_reg_0[4214]),.o(intermediate_reg_1[2107])); 
mux_module mux_module_inst_1_2733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4213]),.i2(intermediate_reg_0[4212]),.o(intermediate_reg_1[2106]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4211]),.i2(intermediate_reg_0[4210]),.o(intermediate_reg_1[2105]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4209]),.i2(intermediate_reg_0[4208]),.o(intermediate_reg_1[2104]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4207]),.i2(intermediate_reg_0[4206]),.o(intermediate_reg_1[2103])); 
fsm fsm_inst_1_2737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4205]),.i2(intermediate_reg_0[4204]),.o(intermediate_reg_1[2102])); 
mux_module mux_module_inst_1_2738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4203]),.i2(intermediate_reg_0[4202]),.o(intermediate_reg_1[2101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4201]),.i2(intermediate_reg_0[4200]),.o(intermediate_reg_1[2100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4199]),.i2(intermediate_reg_0[4198]),.o(intermediate_reg_1[2099]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4197]),.i2(intermediate_reg_0[4196]),.o(intermediate_reg_1[2098])); 
fsm fsm_inst_1_2742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4195]),.i2(intermediate_reg_0[4194]),.o(intermediate_reg_1[2097])); 
mux_module mux_module_inst_1_2743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4193]),.i2(intermediate_reg_0[4192]),.o(intermediate_reg_1[2096]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4191]),.i2(intermediate_reg_0[4190]),.o(intermediate_reg_1[2095])); 
fsm fsm_inst_1_2745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4189]),.i2(intermediate_reg_0[4188]),.o(intermediate_reg_1[2094])); 
mux_module mux_module_inst_1_2746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4187]),.i2(intermediate_reg_0[4186]),.o(intermediate_reg_1[2093]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4185]),.i2(intermediate_reg_0[4184]),.o(intermediate_reg_1[2092]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4183]),.i2(intermediate_reg_0[4182]),.o(intermediate_reg_1[2091])); 
mux_module mux_module_inst_1_2749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4181]),.i2(intermediate_reg_0[4180]),.o(intermediate_reg_1[2090]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4179]),.i2(intermediate_reg_0[4178]),.o(intermediate_reg_1[2089]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4177]),.i2(intermediate_reg_0[4176]),.o(intermediate_reg_1[2088])); 
fsm fsm_inst_1_2752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4175]),.i2(intermediate_reg_0[4174]),.o(intermediate_reg_1[2087])); 
mux_module mux_module_inst_1_2753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4173]),.i2(intermediate_reg_0[4172]),.o(intermediate_reg_1[2086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4171]),.i2(intermediate_reg_0[4170]),.o(intermediate_reg_1[2085]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4169]),.i2(intermediate_reg_0[4168]),.o(intermediate_reg_1[2084])); 
mux_module mux_module_inst_1_2756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4167]),.i2(intermediate_reg_0[4166]),.o(intermediate_reg_1[2083]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4165]),.i2(intermediate_reg_0[4164]),.o(intermediate_reg_1[2082]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4163]),.i2(intermediate_reg_0[4162]),.o(intermediate_reg_1[2081])); 
mux_module mux_module_inst_1_2759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4161]),.i2(intermediate_reg_0[4160]),.o(intermediate_reg_1[2080]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4159]),.i2(intermediate_reg_0[4158]),.o(intermediate_reg_1[2079])); 
mux_module mux_module_inst_1_2761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4157]),.i2(intermediate_reg_0[4156]),.o(intermediate_reg_1[2078]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4155]),.i2(intermediate_reg_0[4154]),.o(intermediate_reg_1[2077]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4153]),.i2(intermediate_reg_0[4152]),.o(intermediate_reg_1[2076])); 
mux_module mux_module_inst_1_2764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4151]),.i2(intermediate_reg_0[4150]),.o(intermediate_reg_1[2075]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4149]),.i2(intermediate_reg_0[4148]),.o(intermediate_reg_1[2074]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4147]),.i2(intermediate_reg_0[4146]),.o(intermediate_reg_1[2073]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4145]),.i2(intermediate_reg_0[4144]),.o(intermediate_reg_1[2072]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4143]),.i2(intermediate_reg_0[4142]),.o(intermediate_reg_1[2071]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4141]),.i2(intermediate_reg_0[4140]),.o(intermediate_reg_1[2070])); 
fsm fsm_inst_1_2770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4139]),.i2(intermediate_reg_0[4138]),.o(intermediate_reg_1[2069])); 
fsm fsm_inst_1_2771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4137]),.i2(intermediate_reg_0[4136]),.o(intermediate_reg_1[2068])); 
fsm fsm_inst_1_2772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4135]),.i2(intermediate_reg_0[4134]),.o(intermediate_reg_1[2067])); 
fsm fsm_inst_1_2773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4133]),.i2(intermediate_reg_0[4132]),.o(intermediate_reg_1[2066])); 
fsm fsm_inst_1_2774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4131]),.i2(intermediate_reg_0[4130]),.o(intermediate_reg_1[2065])); 
mux_module mux_module_inst_1_2775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4129]),.i2(intermediate_reg_0[4128]),.o(intermediate_reg_1[2064]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4127]),.i2(intermediate_reg_0[4126]),.o(intermediate_reg_1[2063]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4125]),.i2(intermediate_reg_0[4124]),.o(intermediate_reg_1[2062]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4123]),.i2(intermediate_reg_0[4122]),.o(intermediate_reg_1[2061])); 
fsm fsm_inst_1_2779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4121]),.i2(intermediate_reg_0[4120]),.o(intermediate_reg_1[2060])); 
fsm fsm_inst_1_2780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4119]),.i2(intermediate_reg_0[4118]),.o(intermediate_reg_1[2059])); 
fsm fsm_inst_1_2781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4117]),.i2(intermediate_reg_0[4116]),.o(intermediate_reg_1[2058])); 
fsm fsm_inst_1_2782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4115]),.i2(intermediate_reg_0[4114]),.o(intermediate_reg_1[2057])); 
mux_module mux_module_inst_1_2783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4113]),.i2(intermediate_reg_0[4112]),.o(intermediate_reg_1[2056]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4111]),.i2(intermediate_reg_0[4110]),.o(intermediate_reg_1[2055]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4109]),.i2(intermediate_reg_0[4108]),.o(intermediate_reg_1[2054])); 
fsm fsm_inst_1_2786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4107]),.i2(intermediate_reg_0[4106]),.o(intermediate_reg_1[2053])); 
mux_module mux_module_inst_1_2787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4105]),.i2(intermediate_reg_0[4104]),.o(intermediate_reg_1[2052]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4103]),.i2(intermediate_reg_0[4102]),.o(intermediate_reg_1[2051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4101]),.i2(intermediate_reg_0[4100]),.o(intermediate_reg_1[2050]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4099]),.i2(intermediate_reg_0[4098]),.o(intermediate_reg_1[2049]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4097]),.i2(intermediate_reg_0[4096]),.o(intermediate_reg_1[2048]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4095]),.i2(intermediate_reg_0[4094]),.o(intermediate_reg_1[2047])); 
fsm fsm_inst_1_2793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4093]),.i2(intermediate_reg_0[4092]),.o(intermediate_reg_1[2046])); 
fsm fsm_inst_1_2794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4091]),.i2(intermediate_reg_0[4090]),.o(intermediate_reg_1[2045])); 
mux_module mux_module_inst_1_2795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4089]),.i2(intermediate_reg_0[4088]),.o(intermediate_reg_1[2044]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4087]),.i2(intermediate_reg_0[4086]),.o(intermediate_reg_1[2043]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4085]),.i2(intermediate_reg_0[4084]),.o(intermediate_reg_1[2042])); 
fsm fsm_inst_1_2798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4083]),.i2(intermediate_reg_0[4082]),.o(intermediate_reg_1[2041])); 
mux_module mux_module_inst_1_2799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4081]),.i2(intermediate_reg_0[4080]),.o(intermediate_reg_1[2040]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4079]),.i2(intermediate_reg_0[4078]),.o(intermediate_reg_1[2039]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4077]),.i2(intermediate_reg_0[4076]),.o(intermediate_reg_1[2038]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4075]),.i2(intermediate_reg_0[4074]),.o(intermediate_reg_1[2037])); 
fsm fsm_inst_1_2803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4073]),.i2(intermediate_reg_0[4072]),.o(intermediate_reg_1[2036])); 
mux_module mux_module_inst_1_2804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4071]),.i2(intermediate_reg_0[4070]),.o(intermediate_reg_1[2035]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4069]),.i2(intermediate_reg_0[4068]),.o(intermediate_reg_1[2034]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4067]),.i2(intermediate_reg_0[4066]),.o(intermediate_reg_1[2033])); 
mux_module mux_module_inst_1_2807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4065]),.i2(intermediate_reg_0[4064]),.o(intermediate_reg_1[2032]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4063]),.i2(intermediate_reg_0[4062]),.o(intermediate_reg_1[2031])); 
fsm fsm_inst_1_2809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4061]),.i2(intermediate_reg_0[4060]),.o(intermediate_reg_1[2030])); 
mux_module mux_module_inst_1_2810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4059]),.i2(intermediate_reg_0[4058]),.o(intermediate_reg_1[2029]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4057]),.i2(intermediate_reg_0[4056]),.o(intermediate_reg_1[2028]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4055]),.i2(intermediate_reg_0[4054]),.o(intermediate_reg_1[2027]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4053]),.i2(intermediate_reg_0[4052]),.o(intermediate_reg_1[2026]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4051]),.i2(intermediate_reg_0[4050]),.o(intermediate_reg_1[2025])); 
fsm fsm_inst_1_2815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4049]),.i2(intermediate_reg_0[4048]),.o(intermediate_reg_1[2024])); 
mux_module mux_module_inst_1_2816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4047]),.i2(intermediate_reg_0[4046]),.o(intermediate_reg_1[2023]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4045]),.i2(intermediate_reg_0[4044]),.o(intermediate_reg_1[2022])); 
mux_module mux_module_inst_1_2818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4043]),.i2(intermediate_reg_0[4042]),.o(intermediate_reg_1[2021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4041]),.i2(intermediate_reg_0[4040]),.o(intermediate_reg_1[2020]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4039]),.i2(intermediate_reg_0[4038]),.o(intermediate_reg_1[2019])); 
fsm fsm_inst_1_2821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4037]),.i2(intermediate_reg_0[4036]),.o(intermediate_reg_1[2018])); 
mux_module mux_module_inst_1_2822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4035]),.i2(intermediate_reg_0[4034]),.o(intermediate_reg_1[2017]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4033]),.i2(intermediate_reg_0[4032]),.o(intermediate_reg_1[2016])); 
mux_module mux_module_inst_1_2824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4031]),.i2(intermediate_reg_0[4030]),.o(intermediate_reg_1[2015]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4029]),.i2(intermediate_reg_0[4028]),.o(intermediate_reg_1[2014]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4027]),.i2(intermediate_reg_0[4026]),.o(intermediate_reg_1[2013]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4025]),.i2(intermediate_reg_0[4024]),.o(intermediate_reg_1[2012]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4023]),.i2(intermediate_reg_0[4022]),.o(intermediate_reg_1[2011])); 
mux_module mux_module_inst_1_2829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4021]),.i2(intermediate_reg_0[4020]),.o(intermediate_reg_1[2010]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4019]),.i2(intermediate_reg_0[4018]),.o(intermediate_reg_1[2009]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4017]),.i2(intermediate_reg_0[4016]),.o(intermediate_reg_1[2008])); 
mux_module mux_module_inst_1_2832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4015]),.i2(intermediate_reg_0[4014]),.o(intermediate_reg_1[2007]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4013]),.i2(intermediate_reg_0[4012]),.o(intermediate_reg_1[2006]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4011]),.i2(intermediate_reg_0[4010]),.o(intermediate_reg_1[2005])); 
mux_module mux_module_inst_1_2835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4009]),.i2(intermediate_reg_0[4008]),.o(intermediate_reg_1[2004]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4007]),.i2(intermediate_reg_0[4006]),.o(intermediate_reg_1[2003])); 
fsm fsm_inst_1_2837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4005]),.i2(intermediate_reg_0[4004]),.o(intermediate_reg_1[2002])); 
fsm fsm_inst_1_2838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4003]),.i2(intermediate_reg_0[4002]),.o(intermediate_reg_1[2001])); 
fsm fsm_inst_1_2839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4001]),.i2(intermediate_reg_0[4000]),.o(intermediate_reg_1[2000])); 
mux_module mux_module_inst_1_2840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3999]),.i2(intermediate_reg_0[3998]),.o(intermediate_reg_1[1999]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3997]),.i2(intermediate_reg_0[3996]),.o(intermediate_reg_1[1998])); 
fsm fsm_inst_1_2842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3995]),.i2(intermediate_reg_0[3994]),.o(intermediate_reg_1[1997])); 
mux_module mux_module_inst_1_2843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3993]),.i2(intermediate_reg_0[3992]),.o(intermediate_reg_1[1996]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3991]),.i2(intermediate_reg_0[3990]),.o(intermediate_reg_1[1995])); 
fsm fsm_inst_1_2845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3989]),.i2(intermediate_reg_0[3988]),.o(intermediate_reg_1[1994])); 
mux_module mux_module_inst_1_2846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3987]),.i2(intermediate_reg_0[3986]),.o(intermediate_reg_1[1993]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3985]),.i2(intermediate_reg_0[3984]),.o(intermediate_reg_1[1992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3983]),.i2(intermediate_reg_0[3982]),.o(intermediate_reg_1[1991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3981]),.i2(intermediate_reg_0[3980]),.o(intermediate_reg_1[1990]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3979]),.i2(intermediate_reg_0[3978]),.o(intermediate_reg_1[1989])); 
fsm fsm_inst_1_2851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3977]),.i2(intermediate_reg_0[3976]),.o(intermediate_reg_1[1988])); 
fsm fsm_inst_1_2852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3975]),.i2(intermediate_reg_0[3974]),.o(intermediate_reg_1[1987])); 
mux_module mux_module_inst_1_2853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3973]),.i2(intermediate_reg_0[3972]),.o(intermediate_reg_1[1986]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3971]),.i2(intermediate_reg_0[3970]),.o(intermediate_reg_1[1985]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3969]),.i2(intermediate_reg_0[3968]),.o(intermediate_reg_1[1984]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3967]),.i2(intermediate_reg_0[3966]),.o(intermediate_reg_1[1983]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3965]),.i2(intermediate_reg_0[3964]),.o(intermediate_reg_1[1982])); 
mux_module mux_module_inst_1_2858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3963]),.i2(intermediate_reg_0[3962]),.o(intermediate_reg_1[1981]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3961]),.i2(intermediate_reg_0[3960]),.o(intermediate_reg_1[1980])); 
fsm fsm_inst_1_2860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3959]),.i2(intermediate_reg_0[3958]),.o(intermediate_reg_1[1979])); 
mux_module mux_module_inst_1_2861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3957]),.i2(intermediate_reg_0[3956]),.o(intermediate_reg_1[1978]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3955]),.i2(intermediate_reg_0[3954]),.o(intermediate_reg_1[1977]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3953]),.i2(intermediate_reg_0[3952]),.o(intermediate_reg_1[1976])); 
mux_module mux_module_inst_1_2864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3951]),.i2(intermediate_reg_0[3950]),.o(intermediate_reg_1[1975]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3949]),.i2(intermediate_reg_0[3948]),.o(intermediate_reg_1[1974])); 
mux_module mux_module_inst_1_2866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3947]),.i2(intermediate_reg_0[3946]),.o(intermediate_reg_1[1973]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3945]),.i2(intermediate_reg_0[3944]),.o(intermediate_reg_1[1972]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3943]),.i2(intermediate_reg_0[3942]),.o(intermediate_reg_1[1971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3941]),.i2(intermediate_reg_0[3940]),.o(intermediate_reg_1[1970]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3939]),.i2(intermediate_reg_0[3938]),.o(intermediate_reg_1[1969])); 
mux_module mux_module_inst_1_2871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3937]),.i2(intermediate_reg_0[3936]),.o(intermediate_reg_1[1968]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3935]),.i2(intermediate_reg_0[3934]),.o(intermediate_reg_1[1967])); 
fsm fsm_inst_1_2873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3933]),.i2(intermediate_reg_0[3932]),.o(intermediate_reg_1[1966])); 
mux_module mux_module_inst_1_2874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3931]),.i2(intermediate_reg_0[3930]),.o(intermediate_reg_1[1965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3929]),.i2(intermediate_reg_0[3928]),.o(intermediate_reg_1[1964]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3927]),.i2(intermediate_reg_0[3926]),.o(intermediate_reg_1[1963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3925]),.i2(intermediate_reg_0[3924]),.o(intermediate_reg_1[1962]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3923]),.i2(intermediate_reg_0[3922]),.o(intermediate_reg_1[1961])); 
fsm fsm_inst_1_2879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3921]),.i2(intermediate_reg_0[3920]),.o(intermediate_reg_1[1960])); 
fsm fsm_inst_1_2880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3919]),.i2(intermediate_reg_0[3918]),.o(intermediate_reg_1[1959])); 
mux_module mux_module_inst_1_2881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3917]),.i2(intermediate_reg_0[3916]),.o(intermediate_reg_1[1958]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3915]),.i2(intermediate_reg_0[3914]),.o(intermediate_reg_1[1957]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3913]),.i2(intermediate_reg_0[3912]),.o(intermediate_reg_1[1956])); 
fsm fsm_inst_1_2884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3911]),.i2(intermediate_reg_0[3910]),.o(intermediate_reg_1[1955])); 
fsm fsm_inst_1_2885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3909]),.i2(intermediate_reg_0[3908]),.o(intermediate_reg_1[1954])); 
mux_module mux_module_inst_1_2886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3907]),.i2(intermediate_reg_0[3906]),.o(intermediate_reg_1[1953]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3905]),.i2(intermediate_reg_0[3904]),.o(intermediate_reg_1[1952]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3903]),.i2(intermediate_reg_0[3902]),.o(intermediate_reg_1[1951]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3901]),.i2(intermediate_reg_0[3900]),.o(intermediate_reg_1[1950])); 
fsm fsm_inst_1_2890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3899]),.i2(intermediate_reg_0[3898]),.o(intermediate_reg_1[1949])); 
mux_module mux_module_inst_1_2891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3897]),.i2(intermediate_reg_0[3896]),.o(intermediate_reg_1[1948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3895]),.i2(intermediate_reg_0[3894]),.o(intermediate_reg_1[1947]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3893]),.i2(intermediate_reg_0[3892]),.o(intermediate_reg_1[1946]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3891]),.i2(intermediate_reg_0[3890]),.o(intermediate_reg_1[1945])); 
mux_module mux_module_inst_1_2895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3889]),.i2(intermediate_reg_0[3888]),.o(intermediate_reg_1[1944]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3887]),.i2(intermediate_reg_0[3886]),.o(intermediate_reg_1[1943]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3885]),.i2(intermediate_reg_0[3884]),.o(intermediate_reg_1[1942])); 
fsm fsm_inst_1_2898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3883]),.i2(intermediate_reg_0[3882]),.o(intermediate_reg_1[1941])); 
fsm fsm_inst_1_2899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3881]),.i2(intermediate_reg_0[3880]),.o(intermediate_reg_1[1940])); 
mux_module mux_module_inst_1_2900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3879]),.i2(intermediate_reg_0[3878]),.o(intermediate_reg_1[1939]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3877]),.i2(intermediate_reg_0[3876]),.o(intermediate_reg_1[1938]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3875]),.i2(intermediate_reg_0[3874]),.o(intermediate_reg_1[1937]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3873]),.i2(intermediate_reg_0[3872]),.o(intermediate_reg_1[1936])); 
mux_module mux_module_inst_1_2904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3871]),.i2(intermediate_reg_0[3870]),.o(intermediate_reg_1[1935]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3869]),.i2(intermediate_reg_0[3868]),.o(intermediate_reg_1[1934]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3867]),.i2(intermediate_reg_0[3866]),.o(intermediate_reg_1[1933])); 
fsm fsm_inst_1_2907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3865]),.i2(intermediate_reg_0[3864]),.o(intermediate_reg_1[1932])); 
fsm fsm_inst_1_2908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3863]),.i2(intermediate_reg_0[3862]),.o(intermediate_reg_1[1931])); 
mux_module mux_module_inst_1_2909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3861]),.i2(intermediate_reg_0[3860]),.o(intermediate_reg_1[1930]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3859]),.i2(intermediate_reg_0[3858]),.o(intermediate_reg_1[1929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3857]),.i2(intermediate_reg_0[3856]),.o(intermediate_reg_1[1928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3855]),.i2(intermediate_reg_0[3854]),.o(intermediate_reg_1[1927]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3853]),.i2(intermediate_reg_0[3852]),.o(intermediate_reg_1[1926]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3851]),.i2(intermediate_reg_0[3850]),.o(intermediate_reg_1[1925])); 
mux_module mux_module_inst_1_2915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3849]),.i2(intermediate_reg_0[3848]),.o(intermediate_reg_1[1924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3847]),.i2(intermediate_reg_0[3846]),.o(intermediate_reg_1[1923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3845]),.i2(intermediate_reg_0[3844]),.o(intermediate_reg_1[1922]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3843]),.i2(intermediate_reg_0[3842]),.o(intermediate_reg_1[1921])); 
fsm fsm_inst_1_2919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3841]),.i2(intermediate_reg_0[3840]),.o(intermediate_reg_1[1920])); 
mux_module mux_module_inst_1_2920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3839]),.i2(intermediate_reg_0[3838]),.o(intermediate_reg_1[1919]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3837]),.i2(intermediate_reg_0[3836]),.o(intermediate_reg_1[1918])); 
mux_module mux_module_inst_1_2922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3835]),.i2(intermediate_reg_0[3834]),.o(intermediate_reg_1[1917]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3833]),.i2(intermediate_reg_0[3832]),.o(intermediate_reg_1[1916]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3831]),.i2(intermediate_reg_0[3830]),.o(intermediate_reg_1[1915])); 
mux_module mux_module_inst_1_2925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3829]),.i2(intermediate_reg_0[3828]),.o(intermediate_reg_1[1914]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3827]),.i2(intermediate_reg_0[3826]),.o(intermediate_reg_1[1913]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3825]),.i2(intermediate_reg_0[3824]),.o(intermediate_reg_1[1912]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3823]),.i2(intermediate_reg_0[3822]),.o(intermediate_reg_1[1911]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3821]),.i2(intermediate_reg_0[3820]),.o(intermediate_reg_1[1910]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3819]),.i2(intermediate_reg_0[3818]),.o(intermediate_reg_1[1909])); 
mux_module mux_module_inst_1_2931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3817]),.i2(intermediate_reg_0[3816]),.o(intermediate_reg_1[1908]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3815]),.i2(intermediate_reg_0[3814]),.o(intermediate_reg_1[1907])); 
fsm fsm_inst_1_2933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3813]),.i2(intermediate_reg_0[3812]),.o(intermediate_reg_1[1906])); 
fsm fsm_inst_1_2934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3811]),.i2(intermediate_reg_0[3810]),.o(intermediate_reg_1[1905])); 
fsm fsm_inst_1_2935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3809]),.i2(intermediate_reg_0[3808]),.o(intermediate_reg_1[1904])); 
fsm fsm_inst_1_2936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3807]),.i2(intermediate_reg_0[3806]),.o(intermediate_reg_1[1903])); 
fsm fsm_inst_1_2937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3805]),.i2(intermediate_reg_0[3804]),.o(intermediate_reg_1[1902])); 
mux_module mux_module_inst_1_2938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3803]),.i2(intermediate_reg_0[3802]),.o(intermediate_reg_1[1901]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3801]),.i2(intermediate_reg_0[3800]),.o(intermediate_reg_1[1900])); 
fsm fsm_inst_1_2940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3799]),.i2(intermediate_reg_0[3798]),.o(intermediate_reg_1[1899])); 
mux_module mux_module_inst_1_2941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3797]),.i2(intermediate_reg_0[3796]),.o(intermediate_reg_1[1898]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3795]),.i2(intermediate_reg_0[3794]),.o(intermediate_reg_1[1897])); 
fsm fsm_inst_1_2943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3793]),.i2(intermediate_reg_0[3792]),.o(intermediate_reg_1[1896])); 
mux_module mux_module_inst_1_2944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3791]),.i2(intermediate_reg_0[3790]),.o(intermediate_reg_1[1895]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3789]),.i2(intermediate_reg_0[3788]),.o(intermediate_reg_1[1894])); 
fsm fsm_inst_1_2946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3787]),.i2(intermediate_reg_0[3786]),.o(intermediate_reg_1[1893])); 
mux_module mux_module_inst_1_2947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3785]),.i2(intermediate_reg_0[3784]),.o(intermediate_reg_1[1892]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3783]),.i2(intermediate_reg_0[3782]),.o(intermediate_reg_1[1891]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3781]),.i2(intermediate_reg_0[3780]),.o(intermediate_reg_1[1890]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3779]),.i2(intermediate_reg_0[3778]),.o(intermediate_reg_1[1889])); 
mux_module mux_module_inst_1_2951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3777]),.i2(intermediate_reg_0[3776]),.o(intermediate_reg_1[1888]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3775]),.i2(intermediate_reg_0[3774]),.o(intermediate_reg_1[1887]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3773]),.i2(intermediate_reg_0[3772]),.o(intermediate_reg_1[1886]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3771]),.i2(intermediate_reg_0[3770]),.o(intermediate_reg_1[1885])); 
fsm fsm_inst_1_2955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3769]),.i2(intermediate_reg_0[3768]),.o(intermediate_reg_1[1884])); 
fsm fsm_inst_1_2956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3767]),.i2(intermediate_reg_0[3766]),.o(intermediate_reg_1[1883])); 
mux_module mux_module_inst_1_2957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3765]),.i2(intermediate_reg_0[3764]),.o(intermediate_reg_1[1882]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3763]),.i2(intermediate_reg_0[3762]),.o(intermediate_reg_1[1881])); 
fsm fsm_inst_1_2959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3761]),.i2(intermediate_reg_0[3760]),.o(intermediate_reg_1[1880])); 
mux_module mux_module_inst_1_2960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3759]),.i2(intermediate_reg_0[3758]),.o(intermediate_reg_1[1879]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3757]),.i2(intermediate_reg_0[3756]),.o(intermediate_reg_1[1878]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3755]),.i2(intermediate_reg_0[3754]),.o(intermediate_reg_1[1877])); 
fsm fsm_inst_1_2963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3753]),.i2(intermediate_reg_0[3752]),.o(intermediate_reg_1[1876])); 
fsm fsm_inst_1_2964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3751]),.i2(intermediate_reg_0[3750]),.o(intermediate_reg_1[1875])); 
mux_module mux_module_inst_1_2965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3749]),.i2(intermediate_reg_0[3748]),.o(intermediate_reg_1[1874]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3747]),.i2(intermediate_reg_0[3746]),.o(intermediate_reg_1[1873])); 
mux_module mux_module_inst_1_2967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3745]),.i2(intermediate_reg_0[3744]),.o(intermediate_reg_1[1872]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3743]),.i2(intermediate_reg_0[3742]),.o(intermediate_reg_1[1871]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3741]),.i2(intermediate_reg_0[3740]),.o(intermediate_reg_1[1870])); 
mux_module mux_module_inst_1_2970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3739]),.i2(intermediate_reg_0[3738]),.o(intermediate_reg_1[1869]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3737]),.i2(intermediate_reg_0[3736]),.o(intermediate_reg_1[1868])); 
mux_module mux_module_inst_1_2972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3735]),.i2(intermediate_reg_0[3734]),.o(intermediate_reg_1[1867]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3733]),.i2(intermediate_reg_0[3732]),.o(intermediate_reg_1[1866])); 
mux_module mux_module_inst_1_2974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3731]),.i2(intermediate_reg_0[3730]),.o(intermediate_reg_1[1865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3729]),.i2(intermediate_reg_0[3728]),.o(intermediate_reg_1[1864]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3727]),.i2(intermediate_reg_0[3726]),.o(intermediate_reg_1[1863]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3725]),.i2(intermediate_reg_0[3724]),.o(intermediate_reg_1[1862]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3723]),.i2(intermediate_reg_0[3722]),.o(intermediate_reg_1[1861])); 
fsm fsm_inst_1_2979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3721]),.i2(intermediate_reg_0[3720]),.o(intermediate_reg_1[1860])); 
fsm fsm_inst_1_2980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3719]),.i2(intermediate_reg_0[3718]),.o(intermediate_reg_1[1859])); 
fsm fsm_inst_1_2981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3717]),.i2(intermediate_reg_0[3716]),.o(intermediate_reg_1[1858])); 
fsm fsm_inst_1_2982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3715]),.i2(intermediate_reg_0[3714]),.o(intermediate_reg_1[1857])); 
mux_module mux_module_inst_1_2983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3713]),.i2(intermediate_reg_0[3712]),.o(intermediate_reg_1[1856]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3711]),.i2(intermediate_reg_0[3710]),.o(intermediate_reg_1[1855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3709]),.i2(intermediate_reg_0[3708]),.o(intermediate_reg_1[1854]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3707]),.i2(intermediate_reg_0[3706]),.o(intermediate_reg_1[1853]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3705]),.i2(intermediate_reg_0[3704]),.o(intermediate_reg_1[1852])); 
mux_module mux_module_inst_1_2988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3703]),.i2(intermediate_reg_0[3702]),.o(intermediate_reg_1[1851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3701]),.i2(intermediate_reg_0[3700]),.o(intermediate_reg_1[1850]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3699]),.i2(intermediate_reg_0[3698]),.o(intermediate_reg_1[1849])); 
fsm fsm_inst_1_2991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3697]),.i2(intermediate_reg_0[3696]),.o(intermediate_reg_1[1848])); 
fsm fsm_inst_1_2992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3695]),.i2(intermediate_reg_0[3694]),.o(intermediate_reg_1[1847])); 
fsm fsm_inst_1_2993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3693]),.i2(intermediate_reg_0[3692]),.o(intermediate_reg_1[1846])); 
fsm fsm_inst_1_2994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3691]),.i2(intermediate_reg_0[3690]),.o(intermediate_reg_1[1845])); 
mux_module mux_module_inst_1_2995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3689]),.i2(intermediate_reg_0[3688]),.o(intermediate_reg_1[1844]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3687]),.i2(intermediate_reg_0[3686]),.o(intermediate_reg_1[1843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3685]),.i2(intermediate_reg_0[3684]),.o(intermediate_reg_1[1842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3683]),.i2(intermediate_reg_0[3682]),.o(intermediate_reg_1[1841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3681]),.i2(intermediate_reg_0[3680]),.o(intermediate_reg_1[1840]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3679]),.i2(intermediate_reg_0[3678]),.o(intermediate_reg_1[1839])); 
mux_module mux_module_inst_1_3001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3677]),.i2(intermediate_reg_0[3676]),.o(intermediate_reg_1[1838]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3675]),.i2(intermediate_reg_0[3674]),.o(intermediate_reg_1[1837]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3673]),.i2(intermediate_reg_0[3672]),.o(intermediate_reg_1[1836]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3671]),.i2(intermediate_reg_0[3670]),.o(intermediate_reg_1[1835]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3669]),.i2(intermediate_reg_0[3668]),.o(intermediate_reg_1[1834]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3667]),.i2(intermediate_reg_0[3666]),.o(intermediate_reg_1[1833])); 
fsm fsm_inst_1_3007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3665]),.i2(intermediate_reg_0[3664]),.o(intermediate_reg_1[1832])); 
fsm fsm_inst_1_3008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3663]),.i2(intermediate_reg_0[3662]),.o(intermediate_reg_1[1831])); 
mux_module mux_module_inst_1_3009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3661]),.i2(intermediate_reg_0[3660]),.o(intermediate_reg_1[1830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3659]),.i2(intermediate_reg_0[3658]),.o(intermediate_reg_1[1829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3657]),.i2(intermediate_reg_0[3656]),.o(intermediate_reg_1[1828]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3655]),.i2(intermediate_reg_0[3654]),.o(intermediate_reg_1[1827]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3653]),.i2(intermediate_reg_0[3652]),.o(intermediate_reg_1[1826]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3651]),.i2(intermediate_reg_0[3650]),.o(intermediate_reg_1[1825]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3649]),.i2(intermediate_reg_0[3648]),.o(intermediate_reg_1[1824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3647]),.i2(intermediate_reg_0[3646]),.o(intermediate_reg_1[1823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3645]),.i2(intermediate_reg_0[3644]),.o(intermediate_reg_1[1822]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3643]),.i2(intermediate_reg_0[3642]),.o(intermediate_reg_1[1821])); 
fsm fsm_inst_1_3019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3641]),.i2(intermediate_reg_0[3640]),.o(intermediate_reg_1[1820])); 
fsm fsm_inst_1_3020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3639]),.i2(intermediate_reg_0[3638]),.o(intermediate_reg_1[1819])); 
mux_module mux_module_inst_1_3021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3637]),.i2(intermediate_reg_0[3636]),.o(intermediate_reg_1[1818]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3635]),.i2(intermediate_reg_0[3634]),.o(intermediate_reg_1[1817]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3633]),.i2(intermediate_reg_0[3632]),.o(intermediate_reg_1[1816]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3631]),.i2(intermediate_reg_0[3630]),.o(intermediate_reg_1[1815])); 
fsm fsm_inst_1_3025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3629]),.i2(intermediate_reg_0[3628]),.o(intermediate_reg_1[1814])); 
mux_module mux_module_inst_1_3026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3627]),.i2(intermediate_reg_0[3626]),.o(intermediate_reg_1[1813]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3625]),.i2(intermediate_reg_0[3624]),.o(intermediate_reg_1[1812])); 
fsm fsm_inst_1_3028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3623]),.i2(intermediate_reg_0[3622]),.o(intermediate_reg_1[1811])); 
mux_module mux_module_inst_1_3029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3621]),.i2(intermediate_reg_0[3620]),.o(intermediate_reg_1[1810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3619]),.i2(intermediate_reg_0[3618]),.o(intermediate_reg_1[1809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3617]),.i2(intermediate_reg_0[3616]),.o(intermediate_reg_1[1808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3615]),.i2(intermediate_reg_0[3614]),.o(intermediate_reg_1[1807]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3613]),.i2(intermediate_reg_0[3612]),.o(intermediate_reg_1[1806]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3611]),.i2(intermediate_reg_0[3610]),.o(intermediate_reg_1[1805])); 
mux_module mux_module_inst_1_3035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3609]),.i2(intermediate_reg_0[3608]),.o(intermediate_reg_1[1804]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3607]),.i2(intermediate_reg_0[3606]),.o(intermediate_reg_1[1803])); 
mux_module mux_module_inst_1_3037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3605]),.i2(intermediate_reg_0[3604]),.o(intermediate_reg_1[1802]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3603]),.i2(intermediate_reg_0[3602]),.o(intermediate_reg_1[1801])); 
fsm fsm_inst_1_3039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3601]),.i2(intermediate_reg_0[3600]),.o(intermediate_reg_1[1800])); 
fsm fsm_inst_1_3040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3599]),.i2(intermediate_reg_0[3598]),.o(intermediate_reg_1[1799])); 
mux_module mux_module_inst_1_3041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3597]),.i2(intermediate_reg_0[3596]),.o(intermediate_reg_1[1798]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3595]),.i2(intermediate_reg_0[3594]),.o(intermediate_reg_1[1797])); 
mux_module mux_module_inst_1_3043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3593]),.i2(intermediate_reg_0[3592]),.o(intermediate_reg_1[1796]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3591]),.i2(intermediate_reg_0[3590]),.o(intermediate_reg_1[1795])); 
mux_module mux_module_inst_1_3045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3589]),.i2(intermediate_reg_0[3588]),.o(intermediate_reg_1[1794]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3587]),.i2(intermediate_reg_0[3586]),.o(intermediate_reg_1[1793])); 
fsm fsm_inst_1_3047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3585]),.i2(intermediate_reg_0[3584]),.o(intermediate_reg_1[1792])); 
fsm fsm_inst_1_3048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3583]),.i2(intermediate_reg_0[3582]),.o(intermediate_reg_1[1791])); 
mux_module mux_module_inst_1_3049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3581]),.i2(intermediate_reg_0[3580]),.o(intermediate_reg_1[1790]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3579]),.i2(intermediate_reg_0[3578]),.o(intermediate_reg_1[1789])); 
fsm fsm_inst_1_3051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3577]),.i2(intermediate_reg_0[3576]),.o(intermediate_reg_1[1788])); 
mux_module mux_module_inst_1_3052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3575]),.i2(intermediate_reg_0[3574]),.o(intermediate_reg_1[1787]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3573]),.i2(intermediate_reg_0[3572]),.o(intermediate_reg_1[1786]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3571]),.i2(intermediate_reg_0[3570]),.o(intermediate_reg_1[1785])); 
fsm fsm_inst_1_3055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3569]),.i2(intermediate_reg_0[3568]),.o(intermediate_reg_1[1784])); 
mux_module mux_module_inst_1_3056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3567]),.i2(intermediate_reg_0[3566]),.o(intermediate_reg_1[1783]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3565]),.i2(intermediate_reg_0[3564]),.o(intermediate_reg_1[1782])); 
fsm fsm_inst_1_3058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3563]),.i2(intermediate_reg_0[3562]),.o(intermediate_reg_1[1781])); 
mux_module mux_module_inst_1_3059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3561]),.i2(intermediate_reg_0[3560]),.o(intermediate_reg_1[1780]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3559]),.i2(intermediate_reg_0[3558]),.o(intermediate_reg_1[1779]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3557]),.i2(intermediate_reg_0[3556]),.o(intermediate_reg_1[1778]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3555]),.i2(intermediate_reg_0[3554]),.o(intermediate_reg_1[1777])); 
fsm fsm_inst_1_3063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3553]),.i2(intermediate_reg_0[3552]),.o(intermediate_reg_1[1776])); 
fsm fsm_inst_1_3064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3551]),.i2(intermediate_reg_0[3550]),.o(intermediate_reg_1[1775])); 
fsm fsm_inst_1_3065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3549]),.i2(intermediate_reg_0[3548]),.o(intermediate_reg_1[1774])); 
fsm fsm_inst_1_3066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3547]),.i2(intermediate_reg_0[3546]),.o(intermediate_reg_1[1773])); 
mux_module mux_module_inst_1_3067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3545]),.i2(intermediate_reg_0[3544]),.o(intermediate_reg_1[1772]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3543]),.i2(intermediate_reg_0[3542]),.o(intermediate_reg_1[1771]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3541]),.i2(intermediate_reg_0[3540]),.o(intermediate_reg_1[1770]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3539]),.i2(intermediate_reg_0[3538]),.o(intermediate_reg_1[1769]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3537]),.i2(intermediate_reg_0[3536]),.o(intermediate_reg_1[1768])); 
mux_module mux_module_inst_1_3072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3535]),.i2(intermediate_reg_0[3534]),.o(intermediate_reg_1[1767]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3533]),.i2(intermediate_reg_0[3532]),.o(intermediate_reg_1[1766]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3531]),.i2(intermediate_reg_0[3530]),.o(intermediate_reg_1[1765])); 
fsm fsm_inst_1_3075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3529]),.i2(intermediate_reg_0[3528]),.o(intermediate_reg_1[1764])); 
mux_module mux_module_inst_1_3076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3527]),.i2(intermediate_reg_0[3526]),.o(intermediate_reg_1[1763]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3525]),.i2(intermediate_reg_0[3524]),.o(intermediate_reg_1[1762])); 
fsm fsm_inst_1_3078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3523]),.i2(intermediate_reg_0[3522]),.o(intermediate_reg_1[1761])); 
fsm fsm_inst_1_3079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3521]),.i2(intermediate_reg_0[3520]),.o(intermediate_reg_1[1760])); 
fsm fsm_inst_1_3080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3519]),.i2(intermediate_reg_0[3518]),.o(intermediate_reg_1[1759])); 
mux_module mux_module_inst_1_3081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3517]),.i2(intermediate_reg_0[3516]),.o(intermediate_reg_1[1758]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3515]),.i2(intermediate_reg_0[3514]),.o(intermediate_reg_1[1757])); 
mux_module mux_module_inst_1_3083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3513]),.i2(intermediate_reg_0[3512]),.o(intermediate_reg_1[1756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3511]),.i2(intermediate_reg_0[3510]),.o(intermediate_reg_1[1755]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3509]),.i2(intermediate_reg_0[3508]),.o(intermediate_reg_1[1754])); 
mux_module mux_module_inst_1_3086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3507]),.i2(intermediate_reg_0[3506]),.o(intermediate_reg_1[1753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3505]),.i2(intermediate_reg_0[3504]),.o(intermediate_reg_1[1752]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3503]),.i2(intermediate_reg_0[3502]),.o(intermediate_reg_1[1751])); 
mux_module mux_module_inst_1_3089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3501]),.i2(intermediate_reg_0[3500]),.o(intermediate_reg_1[1750]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3499]),.i2(intermediate_reg_0[3498]),.o(intermediate_reg_1[1749]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3497]),.i2(intermediate_reg_0[3496]),.o(intermediate_reg_1[1748])); 
fsm fsm_inst_1_3092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3495]),.i2(intermediate_reg_0[3494]),.o(intermediate_reg_1[1747])); 
fsm fsm_inst_1_3093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3493]),.i2(intermediate_reg_0[3492]),.o(intermediate_reg_1[1746])); 
mux_module mux_module_inst_1_3094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3491]),.i2(intermediate_reg_0[3490]),.o(intermediate_reg_1[1745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3489]),.i2(intermediate_reg_0[3488]),.o(intermediate_reg_1[1744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3487]),.i2(intermediate_reg_0[3486]),.o(intermediate_reg_1[1743]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3485]),.i2(intermediate_reg_0[3484]),.o(intermediate_reg_1[1742])); 
fsm fsm_inst_1_3098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3483]),.i2(intermediate_reg_0[3482]),.o(intermediate_reg_1[1741])); 
mux_module mux_module_inst_1_3099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3481]),.i2(intermediate_reg_0[3480]),.o(intermediate_reg_1[1740]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3479]),.i2(intermediate_reg_0[3478]),.o(intermediate_reg_1[1739])); 
mux_module mux_module_inst_1_3101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3477]),.i2(intermediate_reg_0[3476]),.o(intermediate_reg_1[1738]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3475]),.i2(intermediate_reg_0[3474]),.o(intermediate_reg_1[1737])); 
fsm fsm_inst_1_3103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3473]),.i2(intermediate_reg_0[3472]),.o(intermediate_reg_1[1736])); 
mux_module mux_module_inst_1_3104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3471]),.i2(intermediate_reg_0[3470]),.o(intermediate_reg_1[1735]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3469]),.i2(intermediate_reg_0[3468]),.o(intermediate_reg_1[1734]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3467]),.i2(intermediate_reg_0[3466]),.o(intermediate_reg_1[1733])); 
mux_module mux_module_inst_1_3107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3465]),.i2(intermediate_reg_0[3464]),.o(intermediate_reg_1[1732]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3463]),.i2(intermediate_reg_0[3462]),.o(intermediate_reg_1[1731])); 
fsm fsm_inst_1_3109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3461]),.i2(intermediate_reg_0[3460]),.o(intermediate_reg_1[1730])); 
mux_module mux_module_inst_1_3110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3459]),.i2(intermediate_reg_0[3458]),.o(intermediate_reg_1[1729]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3457]),.i2(intermediate_reg_0[3456]),.o(intermediate_reg_1[1728])); 
fsm fsm_inst_1_3112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3455]),.i2(intermediate_reg_0[3454]),.o(intermediate_reg_1[1727])); 
fsm fsm_inst_1_3113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3453]),.i2(intermediate_reg_0[3452]),.o(intermediate_reg_1[1726])); 
fsm fsm_inst_1_3114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3451]),.i2(intermediate_reg_0[3450]),.o(intermediate_reg_1[1725])); 
fsm fsm_inst_1_3115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3449]),.i2(intermediate_reg_0[3448]),.o(intermediate_reg_1[1724])); 
mux_module mux_module_inst_1_3116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3447]),.i2(intermediate_reg_0[3446]),.o(intermediate_reg_1[1723]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3445]),.i2(intermediate_reg_0[3444]),.o(intermediate_reg_1[1722])); 
mux_module mux_module_inst_1_3118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3443]),.i2(intermediate_reg_0[3442]),.o(intermediate_reg_1[1721]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3441]),.i2(intermediate_reg_0[3440]),.o(intermediate_reg_1[1720]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3439]),.i2(intermediate_reg_0[3438]),.o(intermediate_reg_1[1719]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3437]),.i2(intermediate_reg_0[3436]),.o(intermediate_reg_1[1718]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3435]),.i2(intermediate_reg_0[3434]),.o(intermediate_reg_1[1717]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3433]),.i2(intermediate_reg_0[3432]),.o(intermediate_reg_1[1716])); 
fsm fsm_inst_1_3124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3431]),.i2(intermediate_reg_0[3430]),.o(intermediate_reg_1[1715])); 
fsm fsm_inst_1_3125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3429]),.i2(intermediate_reg_0[3428]),.o(intermediate_reg_1[1714])); 
mux_module mux_module_inst_1_3126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3427]),.i2(intermediate_reg_0[3426]),.o(intermediate_reg_1[1713]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3425]),.i2(intermediate_reg_0[3424]),.o(intermediate_reg_1[1712]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3423]),.i2(intermediate_reg_0[3422]),.o(intermediate_reg_1[1711]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3421]),.i2(intermediate_reg_0[3420]),.o(intermediate_reg_1[1710])); 
mux_module mux_module_inst_1_3130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3419]),.i2(intermediate_reg_0[3418]),.o(intermediate_reg_1[1709]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3417]),.i2(intermediate_reg_0[3416]),.o(intermediate_reg_1[1708]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3415]),.i2(intermediate_reg_0[3414]),.o(intermediate_reg_1[1707])); 
fsm fsm_inst_1_3133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3413]),.i2(intermediate_reg_0[3412]),.o(intermediate_reg_1[1706])); 
fsm fsm_inst_1_3134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3411]),.i2(intermediate_reg_0[3410]),.o(intermediate_reg_1[1705])); 
fsm fsm_inst_1_3135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3409]),.i2(intermediate_reg_0[3408]),.o(intermediate_reg_1[1704])); 
fsm fsm_inst_1_3136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3407]),.i2(intermediate_reg_0[3406]),.o(intermediate_reg_1[1703])); 
fsm fsm_inst_1_3137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3405]),.i2(intermediate_reg_0[3404]),.o(intermediate_reg_1[1702])); 
mux_module mux_module_inst_1_3138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3403]),.i2(intermediate_reg_0[3402]),.o(intermediate_reg_1[1701]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3401]),.i2(intermediate_reg_0[3400]),.o(intermediate_reg_1[1700]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3399]),.i2(intermediate_reg_0[3398]),.o(intermediate_reg_1[1699])); 
fsm fsm_inst_1_3141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3397]),.i2(intermediate_reg_0[3396]),.o(intermediate_reg_1[1698])); 
mux_module mux_module_inst_1_3142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3395]),.i2(intermediate_reg_0[3394]),.o(intermediate_reg_1[1697]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3393]),.i2(intermediate_reg_0[3392]),.o(intermediate_reg_1[1696])); 
fsm fsm_inst_1_3144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3391]),.i2(intermediate_reg_0[3390]),.o(intermediate_reg_1[1695])); 
fsm fsm_inst_1_3145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3389]),.i2(intermediate_reg_0[3388]),.o(intermediate_reg_1[1694])); 
fsm fsm_inst_1_3146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3387]),.i2(intermediate_reg_0[3386]),.o(intermediate_reg_1[1693])); 
fsm fsm_inst_1_3147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3385]),.i2(intermediate_reg_0[3384]),.o(intermediate_reg_1[1692])); 
mux_module mux_module_inst_1_3148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3383]),.i2(intermediate_reg_0[3382]),.o(intermediate_reg_1[1691]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3381]),.i2(intermediate_reg_0[3380]),.o(intermediate_reg_1[1690])); 
mux_module mux_module_inst_1_3150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3379]),.i2(intermediate_reg_0[3378]),.o(intermediate_reg_1[1689]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3377]),.i2(intermediate_reg_0[3376]),.o(intermediate_reg_1[1688]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3375]),.i2(intermediate_reg_0[3374]),.o(intermediate_reg_1[1687])); 
fsm fsm_inst_1_3153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3373]),.i2(intermediate_reg_0[3372]),.o(intermediate_reg_1[1686])); 
mux_module mux_module_inst_1_3154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3371]),.i2(intermediate_reg_0[3370]),.o(intermediate_reg_1[1685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3369]),.i2(intermediate_reg_0[3368]),.o(intermediate_reg_1[1684]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3367]),.i2(intermediate_reg_0[3366]),.o(intermediate_reg_1[1683])); 
fsm fsm_inst_1_3157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3365]),.i2(intermediate_reg_0[3364]),.o(intermediate_reg_1[1682])); 
mux_module mux_module_inst_1_3158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3363]),.i2(intermediate_reg_0[3362]),.o(intermediate_reg_1[1681]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3361]),.i2(intermediate_reg_0[3360]),.o(intermediate_reg_1[1680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3359]),.i2(intermediate_reg_0[3358]),.o(intermediate_reg_1[1679]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3357]),.i2(intermediate_reg_0[3356]),.o(intermediate_reg_1[1678])); 
mux_module mux_module_inst_1_3162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3355]),.i2(intermediate_reg_0[3354]),.o(intermediate_reg_1[1677]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3353]),.i2(intermediate_reg_0[3352]),.o(intermediate_reg_1[1676]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3351]),.i2(intermediate_reg_0[3350]),.o(intermediate_reg_1[1675])); 
fsm fsm_inst_1_3165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3349]),.i2(intermediate_reg_0[3348]),.o(intermediate_reg_1[1674])); 
fsm fsm_inst_1_3166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3347]),.i2(intermediate_reg_0[3346]),.o(intermediate_reg_1[1673])); 
mux_module mux_module_inst_1_3167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3345]),.i2(intermediate_reg_0[3344]),.o(intermediate_reg_1[1672]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3343]),.i2(intermediate_reg_0[3342]),.o(intermediate_reg_1[1671])); 
mux_module mux_module_inst_1_3169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3341]),.i2(intermediate_reg_0[3340]),.o(intermediate_reg_1[1670]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3339]),.i2(intermediate_reg_0[3338]),.o(intermediate_reg_1[1669]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3337]),.i2(intermediate_reg_0[3336]),.o(intermediate_reg_1[1668]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3335]),.i2(intermediate_reg_0[3334]),.o(intermediate_reg_1[1667])); 
fsm fsm_inst_1_3173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3333]),.i2(intermediate_reg_0[3332]),.o(intermediate_reg_1[1666])); 
fsm fsm_inst_1_3174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3331]),.i2(intermediate_reg_0[3330]),.o(intermediate_reg_1[1665])); 
mux_module mux_module_inst_1_3175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3329]),.i2(intermediate_reg_0[3328]),.o(intermediate_reg_1[1664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3327]),.i2(intermediate_reg_0[3326]),.o(intermediate_reg_1[1663]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3325]),.i2(intermediate_reg_0[3324]),.o(intermediate_reg_1[1662]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3323]),.i2(intermediate_reg_0[3322]),.o(intermediate_reg_1[1661]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3321]),.i2(intermediate_reg_0[3320]),.o(intermediate_reg_1[1660])); 
fsm fsm_inst_1_3180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3319]),.i2(intermediate_reg_0[3318]),.o(intermediate_reg_1[1659])); 
fsm fsm_inst_1_3181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3317]),.i2(intermediate_reg_0[3316]),.o(intermediate_reg_1[1658])); 
fsm fsm_inst_1_3182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3315]),.i2(intermediate_reg_0[3314]),.o(intermediate_reg_1[1657])); 
mux_module mux_module_inst_1_3183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3313]),.i2(intermediate_reg_0[3312]),.o(intermediate_reg_1[1656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3311]),.i2(intermediate_reg_0[3310]),.o(intermediate_reg_1[1655]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3309]),.i2(intermediate_reg_0[3308]),.o(intermediate_reg_1[1654]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3307]),.i2(intermediate_reg_0[3306]),.o(intermediate_reg_1[1653])); 
fsm fsm_inst_1_3187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3305]),.i2(intermediate_reg_0[3304]),.o(intermediate_reg_1[1652])); 
fsm fsm_inst_1_3188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3303]),.i2(intermediate_reg_0[3302]),.o(intermediate_reg_1[1651])); 
fsm fsm_inst_1_3189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3301]),.i2(intermediate_reg_0[3300]),.o(intermediate_reg_1[1650])); 
fsm fsm_inst_1_3190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3299]),.i2(intermediate_reg_0[3298]),.o(intermediate_reg_1[1649])); 
mux_module mux_module_inst_1_3191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3297]),.i2(intermediate_reg_0[3296]),.o(intermediate_reg_1[1648]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3295]),.i2(intermediate_reg_0[3294]),.o(intermediate_reg_1[1647]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3293]),.i2(intermediate_reg_0[3292]),.o(intermediate_reg_1[1646])); 
fsm fsm_inst_1_3194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3291]),.i2(intermediate_reg_0[3290]),.o(intermediate_reg_1[1645])); 
mux_module mux_module_inst_1_3195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3289]),.i2(intermediate_reg_0[3288]),.o(intermediate_reg_1[1644]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3287]),.i2(intermediate_reg_0[3286]),.o(intermediate_reg_1[1643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3285]),.i2(intermediate_reg_0[3284]),.o(intermediate_reg_1[1642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3283]),.i2(intermediate_reg_0[3282]),.o(intermediate_reg_1[1641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3281]),.i2(intermediate_reg_0[3280]),.o(intermediate_reg_1[1640]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3279]),.i2(intermediate_reg_0[3278]),.o(intermediate_reg_1[1639])); 
mux_module mux_module_inst_1_3201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3277]),.i2(intermediate_reg_0[3276]),.o(intermediate_reg_1[1638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3275]),.i2(intermediate_reg_0[3274]),.o(intermediate_reg_1[1637])); 
fsm fsm_inst_1_3203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3273]),.i2(intermediate_reg_0[3272]),.o(intermediate_reg_1[1636])); 
mux_module mux_module_inst_1_3204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3271]),.i2(intermediate_reg_0[3270]),.o(intermediate_reg_1[1635]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3269]),.i2(intermediate_reg_0[3268]),.o(intermediate_reg_1[1634]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3267]),.i2(intermediate_reg_0[3266]),.o(intermediate_reg_1[1633])); 
fsm fsm_inst_1_3207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3265]),.i2(intermediate_reg_0[3264]),.o(intermediate_reg_1[1632])); 
mux_module mux_module_inst_1_3208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3263]),.i2(intermediate_reg_0[3262]),.o(intermediate_reg_1[1631]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3261]),.i2(intermediate_reg_0[3260]),.o(intermediate_reg_1[1630])); 
mux_module mux_module_inst_1_3210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3259]),.i2(intermediate_reg_0[3258]),.o(intermediate_reg_1[1629]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3257]),.i2(intermediate_reg_0[3256]),.o(intermediate_reg_1[1628])); 
fsm fsm_inst_1_3212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3255]),.i2(intermediate_reg_0[3254]),.o(intermediate_reg_1[1627])); 
mux_module mux_module_inst_1_3213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3253]),.i2(intermediate_reg_0[3252]),.o(intermediate_reg_1[1626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3251]),.i2(intermediate_reg_0[3250]),.o(intermediate_reg_1[1625])); 
mux_module mux_module_inst_1_3215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3249]),.i2(intermediate_reg_0[3248]),.o(intermediate_reg_1[1624]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3247]),.i2(intermediate_reg_0[3246]),.o(intermediate_reg_1[1623])); 
mux_module mux_module_inst_1_3217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3245]),.i2(intermediate_reg_0[3244]),.o(intermediate_reg_1[1622]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3243]),.i2(intermediate_reg_0[3242]),.o(intermediate_reg_1[1621])); 
fsm fsm_inst_1_3219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3241]),.i2(intermediate_reg_0[3240]),.o(intermediate_reg_1[1620])); 
fsm fsm_inst_1_3220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3239]),.i2(intermediate_reg_0[3238]),.o(intermediate_reg_1[1619])); 
fsm fsm_inst_1_3221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3237]),.i2(intermediate_reg_0[3236]),.o(intermediate_reg_1[1618])); 
fsm fsm_inst_1_3222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3235]),.i2(intermediate_reg_0[3234]),.o(intermediate_reg_1[1617])); 
mux_module mux_module_inst_1_3223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3233]),.i2(intermediate_reg_0[3232]),.o(intermediate_reg_1[1616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3231]),.i2(intermediate_reg_0[3230]),.o(intermediate_reg_1[1615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3229]),.i2(intermediate_reg_0[3228]),.o(intermediate_reg_1[1614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3227]),.i2(intermediate_reg_0[3226]),.o(intermediate_reg_1[1613]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3225]),.i2(intermediate_reg_0[3224]),.o(intermediate_reg_1[1612])); 
fsm fsm_inst_1_3228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3223]),.i2(intermediate_reg_0[3222]),.o(intermediate_reg_1[1611])); 
fsm fsm_inst_1_3229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3221]),.i2(intermediate_reg_0[3220]),.o(intermediate_reg_1[1610])); 
fsm fsm_inst_1_3230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3219]),.i2(intermediate_reg_0[3218]),.o(intermediate_reg_1[1609])); 
mux_module mux_module_inst_1_3231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3217]),.i2(intermediate_reg_0[3216]),.o(intermediate_reg_1[1608]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3215]),.i2(intermediate_reg_0[3214]),.o(intermediate_reg_1[1607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3213]),.i2(intermediate_reg_0[3212]),.o(intermediate_reg_1[1606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3211]),.i2(intermediate_reg_0[3210]),.o(intermediate_reg_1[1605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3209]),.i2(intermediate_reg_0[3208]),.o(intermediate_reg_1[1604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3207]),.i2(intermediate_reg_0[3206]),.o(intermediate_reg_1[1603]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3205]),.i2(intermediate_reg_0[3204]),.o(intermediate_reg_1[1602])); 
fsm fsm_inst_1_3238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3203]),.i2(intermediate_reg_0[3202]),.o(intermediate_reg_1[1601])); 
fsm fsm_inst_1_3239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3201]),.i2(intermediate_reg_0[3200]),.o(intermediate_reg_1[1600])); 
fsm fsm_inst_1_3240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3199]),.i2(intermediate_reg_0[3198]),.o(intermediate_reg_1[1599])); 
fsm fsm_inst_1_3241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3197]),.i2(intermediate_reg_0[3196]),.o(intermediate_reg_1[1598])); 
mux_module mux_module_inst_1_3242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3195]),.i2(intermediate_reg_0[3194]),.o(intermediate_reg_1[1597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3193]),.i2(intermediate_reg_0[3192]),.o(intermediate_reg_1[1596]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3191]),.i2(intermediate_reg_0[3190]),.o(intermediate_reg_1[1595]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3189]),.i2(intermediate_reg_0[3188]),.o(intermediate_reg_1[1594]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3187]),.i2(intermediate_reg_0[3186]),.o(intermediate_reg_1[1593])); 
mux_module mux_module_inst_1_3247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3185]),.i2(intermediate_reg_0[3184]),.o(intermediate_reg_1[1592]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3183]),.i2(intermediate_reg_0[3182]),.o(intermediate_reg_1[1591])); 
fsm fsm_inst_1_3249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3181]),.i2(intermediate_reg_0[3180]),.o(intermediate_reg_1[1590])); 
fsm fsm_inst_1_3250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3179]),.i2(intermediate_reg_0[3178]),.o(intermediate_reg_1[1589])); 
fsm fsm_inst_1_3251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3177]),.i2(intermediate_reg_0[3176]),.o(intermediate_reg_1[1588])); 
fsm fsm_inst_1_3252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3175]),.i2(intermediate_reg_0[3174]),.o(intermediate_reg_1[1587])); 
fsm fsm_inst_1_3253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3173]),.i2(intermediate_reg_0[3172]),.o(intermediate_reg_1[1586])); 
mux_module mux_module_inst_1_3254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3171]),.i2(intermediate_reg_0[3170]),.o(intermediate_reg_1[1585]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3169]),.i2(intermediate_reg_0[3168]),.o(intermediate_reg_1[1584])); 
fsm fsm_inst_1_3256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3167]),.i2(intermediate_reg_0[3166]),.o(intermediate_reg_1[1583])); 
mux_module mux_module_inst_1_3257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3165]),.i2(intermediate_reg_0[3164]),.o(intermediate_reg_1[1582]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3163]),.i2(intermediate_reg_0[3162]),.o(intermediate_reg_1[1581])); 
fsm fsm_inst_1_3259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3161]),.i2(intermediate_reg_0[3160]),.o(intermediate_reg_1[1580])); 
mux_module mux_module_inst_1_3260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3159]),.i2(intermediate_reg_0[3158]),.o(intermediate_reg_1[1579]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3157]),.i2(intermediate_reg_0[3156]),.o(intermediate_reg_1[1578])); 
fsm fsm_inst_1_3262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3155]),.i2(intermediate_reg_0[3154]),.o(intermediate_reg_1[1577])); 
mux_module mux_module_inst_1_3263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3153]),.i2(intermediate_reg_0[3152]),.o(intermediate_reg_1[1576]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3151]),.i2(intermediate_reg_0[3150]),.o(intermediate_reg_1[1575])); 
mux_module mux_module_inst_1_3265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3149]),.i2(intermediate_reg_0[3148]),.o(intermediate_reg_1[1574]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3147]),.i2(intermediate_reg_0[3146]),.o(intermediate_reg_1[1573])); 
mux_module mux_module_inst_1_3267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3145]),.i2(intermediate_reg_0[3144]),.o(intermediate_reg_1[1572]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3143]),.i2(intermediate_reg_0[3142]),.o(intermediate_reg_1[1571]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3141]),.i2(intermediate_reg_0[3140]),.o(intermediate_reg_1[1570]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3139]),.i2(intermediate_reg_0[3138]),.o(intermediate_reg_1[1569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3137]),.i2(intermediate_reg_0[3136]),.o(intermediate_reg_1[1568]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3135]),.i2(intermediate_reg_0[3134]),.o(intermediate_reg_1[1567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3133]),.i2(intermediate_reg_0[3132]),.o(intermediate_reg_1[1566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3131]),.i2(intermediate_reg_0[3130]),.o(intermediate_reg_1[1565]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3129]),.i2(intermediate_reg_0[3128]),.o(intermediate_reg_1[1564])); 
mux_module mux_module_inst_1_3276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3127]),.i2(intermediate_reg_0[3126]),.o(intermediate_reg_1[1563]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3125]),.i2(intermediate_reg_0[3124]),.o(intermediate_reg_1[1562]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3123]),.i2(intermediate_reg_0[3122]),.o(intermediate_reg_1[1561]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3121]),.i2(intermediate_reg_0[3120]),.o(intermediate_reg_1[1560])); 
fsm fsm_inst_1_3280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3119]),.i2(intermediate_reg_0[3118]),.o(intermediate_reg_1[1559])); 
fsm fsm_inst_1_3281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3117]),.i2(intermediate_reg_0[3116]),.o(intermediate_reg_1[1558])); 
mux_module mux_module_inst_1_3282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3115]),.i2(intermediate_reg_0[3114]),.o(intermediate_reg_1[1557]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3113]),.i2(intermediate_reg_0[3112]),.o(intermediate_reg_1[1556]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3111]),.i2(intermediate_reg_0[3110]),.o(intermediate_reg_1[1555]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3109]),.i2(intermediate_reg_0[3108]),.o(intermediate_reg_1[1554])); 
mux_module mux_module_inst_1_3286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3107]),.i2(intermediate_reg_0[3106]),.o(intermediate_reg_1[1553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3105]),.i2(intermediate_reg_0[3104]),.o(intermediate_reg_1[1552]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3103]),.i2(intermediate_reg_0[3102]),.o(intermediate_reg_1[1551])); 
fsm fsm_inst_1_3289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3101]),.i2(intermediate_reg_0[3100]),.o(intermediate_reg_1[1550])); 
mux_module mux_module_inst_1_3290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3099]),.i2(intermediate_reg_0[3098]),.o(intermediate_reg_1[1549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3097]),.i2(intermediate_reg_0[3096]),.o(intermediate_reg_1[1548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3095]),.i2(intermediate_reg_0[3094]),.o(intermediate_reg_1[1547]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3093]),.i2(intermediate_reg_0[3092]),.o(intermediate_reg_1[1546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3091]),.i2(intermediate_reg_0[3090]),.o(intermediate_reg_1[1545]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3089]),.i2(intermediate_reg_0[3088]),.o(intermediate_reg_1[1544])); 
mux_module mux_module_inst_1_3296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3087]),.i2(intermediate_reg_0[3086]),.o(intermediate_reg_1[1543]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3085]),.i2(intermediate_reg_0[3084]),.o(intermediate_reg_1[1542]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3083]),.i2(intermediate_reg_0[3082]),.o(intermediate_reg_1[1541]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3081]),.i2(intermediate_reg_0[3080]),.o(intermediate_reg_1[1540])); 
fsm fsm_inst_1_3300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3079]),.i2(intermediate_reg_0[3078]),.o(intermediate_reg_1[1539])); 
mux_module mux_module_inst_1_3301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3077]),.i2(intermediate_reg_0[3076]),.o(intermediate_reg_1[1538]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3075]),.i2(intermediate_reg_0[3074]),.o(intermediate_reg_1[1537])); 
mux_module mux_module_inst_1_3303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3073]),.i2(intermediate_reg_0[3072]),.o(intermediate_reg_1[1536]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3071]),.i2(intermediate_reg_0[3070]),.o(intermediate_reg_1[1535])); 
mux_module mux_module_inst_1_3305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3069]),.i2(intermediate_reg_0[3068]),.o(intermediate_reg_1[1534]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3067]),.i2(intermediate_reg_0[3066]),.o(intermediate_reg_1[1533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3065]),.i2(intermediate_reg_0[3064]),.o(intermediate_reg_1[1532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3063]),.i2(intermediate_reg_0[3062]),.o(intermediate_reg_1[1531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3061]),.i2(intermediate_reg_0[3060]),.o(intermediate_reg_1[1530]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3059]),.i2(intermediate_reg_0[3058]),.o(intermediate_reg_1[1529])); 
fsm fsm_inst_1_3311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3057]),.i2(intermediate_reg_0[3056]),.o(intermediate_reg_1[1528])); 
mux_module mux_module_inst_1_3312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3055]),.i2(intermediate_reg_0[3054]),.o(intermediate_reg_1[1527]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3053]),.i2(intermediate_reg_0[3052]),.o(intermediate_reg_1[1526])); 
mux_module mux_module_inst_1_3314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3051]),.i2(intermediate_reg_0[3050]),.o(intermediate_reg_1[1525]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3049]),.i2(intermediate_reg_0[3048]),.o(intermediate_reg_1[1524]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3047]),.i2(intermediate_reg_0[3046]),.o(intermediate_reg_1[1523])); 
fsm fsm_inst_1_3317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3045]),.i2(intermediate_reg_0[3044]),.o(intermediate_reg_1[1522])); 
mux_module mux_module_inst_1_3318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3043]),.i2(intermediate_reg_0[3042]),.o(intermediate_reg_1[1521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3041]),.i2(intermediate_reg_0[3040]),.o(intermediate_reg_1[1520]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3039]),.i2(intermediate_reg_0[3038]),.o(intermediate_reg_1[1519])); 
fsm fsm_inst_1_3321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3037]),.i2(intermediate_reg_0[3036]),.o(intermediate_reg_1[1518])); 
fsm fsm_inst_1_3322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3035]),.i2(intermediate_reg_0[3034]),.o(intermediate_reg_1[1517])); 
fsm fsm_inst_1_3323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3033]),.i2(intermediate_reg_0[3032]),.o(intermediate_reg_1[1516])); 
mux_module mux_module_inst_1_3324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3031]),.i2(intermediate_reg_0[3030]),.o(intermediate_reg_1[1515]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3029]),.i2(intermediate_reg_0[3028]),.o(intermediate_reg_1[1514])); 
mux_module mux_module_inst_1_3326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3027]),.i2(intermediate_reg_0[3026]),.o(intermediate_reg_1[1513]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3025]),.i2(intermediate_reg_0[3024]),.o(intermediate_reg_1[1512])); 
fsm fsm_inst_1_3328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3023]),.i2(intermediate_reg_0[3022]),.o(intermediate_reg_1[1511])); 
mux_module mux_module_inst_1_3329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3021]),.i2(intermediate_reg_0[3020]),.o(intermediate_reg_1[1510]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3019]),.i2(intermediate_reg_0[3018]),.o(intermediate_reg_1[1509])); 
fsm fsm_inst_1_3331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3017]),.i2(intermediate_reg_0[3016]),.o(intermediate_reg_1[1508])); 
mux_module mux_module_inst_1_3332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3015]),.i2(intermediate_reg_0[3014]),.o(intermediate_reg_1[1507]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3013]),.i2(intermediate_reg_0[3012]),.o(intermediate_reg_1[1506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3011]),.i2(intermediate_reg_0[3010]),.o(intermediate_reg_1[1505]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3009]),.i2(intermediate_reg_0[3008]),.o(intermediate_reg_1[1504])); 
fsm fsm_inst_1_3336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3007]),.i2(intermediate_reg_0[3006]),.o(intermediate_reg_1[1503])); 
mux_module mux_module_inst_1_3337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3005]),.i2(intermediate_reg_0[3004]),.o(intermediate_reg_1[1502]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3003]),.i2(intermediate_reg_0[3002]),.o(intermediate_reg_1[1501])); 
mux_module mux_module_inst_1_3339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3001]),.i2(intermediate_reg_0[3000]),.o(intermediate_reg_1[1500]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2999]),.i2(intermediate_reg_0[2998]),.o(intermediate_reg_1[1499]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2997]),.i2(intermediate_reg_0[2996]),.o(intermediate_reg_1[1498]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2995]),.i2(intermediate_reg_0[2994]),.o(intermediate_reg_1[1497]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2993]),.i2(intermediate_reg_0[2992]),.o(intermediate_reg_1[1496])); 
fsm fsm_inst_1_3344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2991]),.i2(intermediate_reg_0[2990]),.o(intermediate_reg_1[1495])); 
fsm fsm_inst_1_3345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2989]),.i2(intermediate_reg_0[2988]),.o(intermediate_reg_1[1494])); 
mux_module mux_module_inst_1_3346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2987]),.i2(intermediate_reg_0[2986]),.o(intermediate_reg_1[1493]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2985]),.i2(intermediate_reg_0[2984]),.o(intermediate_reg_1[1492])); 
fsm fsm_inst_1_3348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2983]),.i2(intermediate_reg_0[2982]),.o(intermediate_reg_1[1491])); 
fsm fsm_inst_1_3349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2981]),.i2(intermediate_reg_0[2980]),.o(intermediate_reg_1[1490])); 
fsm fsm_inst_1_3350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2979]),.i2(intermediate_reg_0[2978]),.o(intermediate_reg_1[1489])); 
fsm fsm_inst_1_3351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2977]),.i2(intermediate_reg_0[2976]),.o(intermediate_reg_1[1488])); 
mux_module mux_module_inst_1_3352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2975]),.i2(intermediate_reg_0[2974]),.o(intermediate_reg_1[1487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2973]),.i2(intermediate_reg_0[2972]),.o(intermediate_reg_1[1486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2971]),.i2(intermediate_reg_0[2970]),.o(intermediate_reg_1[1485]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2969]),.i2(intermediate_reg_0[2968]),.o(intermediate_reg_1[1484])); 
mux_module mux_module_inst_1_3356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2967]),.i2(intermediate_reg_0[2966]),.o(intermediate_reg_1[1483]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2965]),.i2(intermediate_reg_0[2964]),.o(intermediate_reg_1[1482])); 
fsm fsm_inst_1_3358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2963]),.i2(intermediate_reg_0[2962]),.o(intermediate_reg_1[1481])); 
mux_module mux_module_inst_1_3359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2961]),.i2(intermediate_reg_0[2960]),.o(intermediate_reg_1[1480]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2959]),.i2(intermediate_reg_0[2958]),.o(intermediate_reg_1[1479])); 
mux_module mux_module_inst_1_3361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2957]),.i2(intermediate_reg_0[2956]),.o(intermediate_reg_1[1478]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2955]),.i2(intermediate_reg_0[2954]),.o(intermediate_reg_1[1477])); 
mux_module mux_module_inst_1_3363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2953]),.i2(intermediate_reg_0[2952]),.o(intermediate_reg_1[1476]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2951]),.i2(intermediate_reg_0[2950]),.o(intermediate_reg_1[1475])); 
mux_module mux_module_inst_1_3365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2949]),.i2(intermediate_reg_0[2948]),.o(intermediate_reg_1[1474]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2947]),.i2(intermediate_reg_0[2946]),.o(intermediate_reg_1[1473])); 
fsm fsm_inst_1_3367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2945]),.i2(intermediate_reg_0[2944]),.o(intermediate_reg_1[1472])); 
mux_module mux_module_inst_1_3368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2943]),.i2(intermediate_reg_0[2942]),.o(intermediate_reg_1[1471]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2941]),.i2(intermediate_reg_0[2940]),.o(intermediate_reg_1[1470])); 
fsm fsm_inst_1_3370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2939]),.i2(intermediate_reg_0[2938]),.o(intermediate_reg_1[1469])); 
fsm fsm_inst_1_3371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2937]),.i2(intermediate_reg_0[2936]),.o(intermediate_reg_1[1468])); 
fsm fsm_inst_1_3372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2935]),.i2(intermediate_reg_0[2934]),.o(intermediate_reg_1[1467])); 
mux_module mux_module_inst_1_3373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2933]),.i2(intermediate_reg_0[2932]),.o(intermediate_reg_1[1466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2931]),.i2(intermediate_reg_0[2930]),.o(intermediate_reg_1[1465]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2929]),.i2(intermediate_reg_0[2928]),.o(intermediate_reg_1[1464]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2927]),.i2(intermediate_reg_0[2926]),.o(intermediate_reg_1[1463])); 
fsm fsm_inst_1_3377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2925]),.i2(intermediate_reg_0[2924]),.o(intermediate_reg_1[1462])); 
mux_module mux_module_inst_1_3378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2923]),.i2(intermediate_reg_0[2922]),.o(intermediate_reg_1[1461]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2921]),.i2(intermediate_reg_0[2920]),.o(intermediate_reg_1[1460])); 
fsm fsm_inst_1_3380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2919]),.i2(intermediate_reg_0[2918]),.o(intermediate_reg_1[1459])); 
mux_module mux_module_inst_1_3381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2917]),.i2(intermediate_reg_0[2916]),.o(intermediate_reg_1[1458]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2915]),.i2(intermediate_reg_0[2914]),.o(intermediate_reg_1[1457])); 
fsm fsm_inst_1_3383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2913]),.i2(intermediate_reg_0[2912]),.o(intermediate_reg_1[1456])); 
fsm fsm_inst_1_3384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2911]),.i2(intermediate_reg_0[2910]),.o(intermediate_reg_1[1455])); 
fsm fsm_inst_1_3385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2909]),.i2(intermediate_reg_0[2908]),.o(intermediate_reg_1[1454])); 
fsm fsm_inst_1_3386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2907]),.i2(intermediate_reg_0[2906]),.o(intermediate_reg_1[1453])); 
fsm fsm_inst_1_3387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2905]),.i2(intermediate_reg_0[2904]),.o(intermediate_reg_1[1452])); 
mux_module mux_module_inst_1_3388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2903]),.i2(intermediate_reg_0[2902]),.o(intermediate_reg_1[1451]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2901]),.i2(intermediate_reg_0[2900]),.o(intermediate_reg_1[1450])); 
fsm fsm_inst_1_3390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2899]),.i2(intermediate_reg_0[2898]),.o(intermediate_reg_1[1449])); 
mux_module mux_module_inst_1_3391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2897]),.i2(intermediate_reg_0[2896]),.o(intermediate_reg_1[1448]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2895]),.i2(intermediate_reg_0[2894]),.o(intermediate_reg_1[1447])); 
fsm fsm_inst_1_3393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2893]),.i2(intermediate_reg_0[2892]),.o(intermediate_reg_1[1446])); 
fsm fsm_inst_1_3394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2891]),.i2(intermediate_reg_0[2890]),.o(intermediate_reg_1[1445])); 
fsm fsm_inst_1_3395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2889]),.i2(intermediate_reg_0[2888]),.o(intermediate_reg_1[1444])); 
fsm fsm_inst_1_3396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2887]),.i2(intermediate_reg_0[2886]),.o(intermediate_reg_1[1443])); 
mux_module mux_module_inst_1_3397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2885]),.i2(intermediate_reg_0[2884]),.o(intermediate_reg_1[1442]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2883]),.i2(intermediate_reg_0[2882]),.o(intermediate_reg_1[1441])); 
fsm fsm_inst_1_3399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2881]),.i2(intermediate_reg_0[2880]),.o(intermediate_reg_1[1440])); 
mux_module mux_module_inst_1_3400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2879]),.i2(intermediate_reg_0[2878]),.o(intermediate_reg_1[1439]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2877]),.i2(intermediate_reg_0[2876]),.o(intermediate_reg_1[1438])); 
fsm fsm_inst_1_3402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2875]),.i2(intermediate_reg_0[2874]),.o(intermediate_reg_1[1437])); 
mux_module mux_module_inst_1_3403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2873]),.i2(intermediate_reg_0[2872]),.o(intermediate_reg_1[1436]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2871]),.i2(intermediate_reg_0[2870]),.o(intermediate_reg_1[1435])); 
mux_module mux_module_inst_1_3405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2869]),.i2(intermediate_reg_0[2868]),.o(intermediate_reg_1[1434]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2867]),.i2(intermediate_reg_0[2866]),.o(intermediate_reg_1[1433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2865]),.i2(intermediate_reg_0[2864]),.o(intermediate_reg_1[1432]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2863]),.i2(intermediate_reg_0[2862]),.o(intermediate_reg_1[1431]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2861]),.i2(intermediate_reg_0[2860]),.o(intermediate_reg_1[1430])); 
fsm fsm_inst_1_3410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2859]),.i2(intermediate_reg_0[2858]),.o(intermediate_reg_1[1429])); 
fsm fsm_inst_1_3411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2857]),.i2(intermediate_reg_0[2856]),.o(intermediate_reg_1[1428])); 
fsm fsm_inst_1_3412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2855]),.i2(intermediate_reg_0[2854]),.o(intermediate_reg_1[1427])); 
mux_module mux_module_inst_1_3413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2853]),.i2(intermediate_reg_0[2852]),.o(intermediate_reg_1[1426]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2851]),.i2(intermediate_reg_0[2850]),.o(intermediate_reg_1[1425])); 
fsm fsm_inst_1_3415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2849]),.i2(intermediate_reg_0[2848]),.o(intermediate_reg_1[1424])); 
mux_module mux_module_inst_1_3416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2847]),.i2(intermediate_reg_0[2846]),.o(intermediate_reg_1[1423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2845]),.i2(intermediate_reg_0[2844]),.o(intermediate_reg_1[1422]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2843]),.i2(intermediate_reg_0[2842]),.o(intermediate_reg_1[1421]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2841]),.i2(intermediate_reg_0[2840]),.o(intermediate_reg_1[1420])); 
fsm fsm_inst_1_3420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2839]),.i2(intermediate_reg_0[2838]),.o(intermediate_reg_1[1419])); 
fsm fsm_inst_1_3421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2837]),.i2(intermediate_reg_0[2836]),.o(intermediate_reg_1[1418])); 
mux_module mux_module_inst_1_3422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2835]),.i2(intermediate_reg_0[2834]),.o(intermediate_reg_1[1417]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2833]),.i2(intermediate_reg_0[2832]),.o(intermediate_reg_1[1416])); 
fsm fsm_inst_1_3424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2831]),.i2(intermediate_reg_0[2830]),.o(intermediate_reg_1[1415])); 
fsm fsm_inst_1_3425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2829]),.i2(intermediate_reg_0[2828]),.o(intermediate_reg_1[1414])); 
fsm fsm_inst_1_3426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2827]),.i2(intermediate_reg_0[2826]),.o(intermediate_reg_1[1413])); 
mux_module mux_module_inst_1_3427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2825]),.i2(intermediate_reg_0[2824]),.o(intermediate_reg_1[1412]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2823]),.i2(intermediate_reg_0[2822]),.o(intermediate_reg_1[1411]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2821]),.i2(intermediate_reg_0[2820]),.o(intermediate_reg_1[1410])); 
fsm fsm_inst_1_3430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2819]),.i2(intermediate_reg_0[2818]),.o(intermediate_reg_1[1409])); 
fsm fsm_inst_1_3431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2817]),.i2(intermediate_reg_0[2816]),.o(intermediate_reg_1[1408])); 
fsm fsm_inst_1_3432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2815]),.i2(intermediate_reg_0[2814]),.o(intermediate_reg_1[1407])); 
mux_module mux_module_inst_1_3433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2813]),.i2(intermediate_reg_0[2812]),.o(intermediate_reg_1[1406]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2811]),.i2(intermediate_reg_0[2810]),.o(intermediate_reg_1[1405])); 
mux_module mux_module_inst_1_3435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2809]),.i2(intermediate_reg_0[2808]),.o(intermediate_reg_1[1404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2807]),.i2(intermediate_reg_0[2806]),.o(intermediate_reg_1[1403])); 
fsm fsm_inst_1_3437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2805]),.i2(intermediate_reg_0[2804]),.o(intermediate_reg_1[1402])); 
fsm fsm_inst_1_3438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2803]),.i2(intermediate_reg_0[2802]),.o(intermediate_reg_1[1401])); 
mux_module mux_module_inst_1_3439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2801]),.i2(intermediate_reg_0[2800]),.o(intermediate_reg_1[1400]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2799]),.i2(intermediate_reg_0[2798]),.o(intermediate_reg_1[1399])); 
fsm fsm_inst_1_3441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2797]),.i2(intermediate_reg_0[2796]),.o(intermediate_reg_1[1398])); 
fsm fsm_inst_1_3442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2795]),.i2(intermediate_reg_0[2794]),.o(intermediate_reg_1[1397])); 
mux_module mux_module_inst_1_3443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2793]),.i2(intermediate_reg_0[2792]),.o(intermediate_reg_1[1396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2791]),.i2(intermediate_reg_0[2790]),.o(intermediate_reg_1[1395]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2789]),.i2(intermediate_reg_0[2788]),.o(intermediate_reg_1[1394])); 
mux_module mux_module_inst_1_3446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2787]),.i2(intermediate_reg_0[2786]),.o(intermediate_reg_1[1393]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2785]),.i2(intermediate_reg_0[2784]),.o(intermediate_reg_1[1392]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2783]),.i2(intermediate_reg_0[2782]),.o(intermediate_reg_1[1391])); 
fsm fsm_inst_1_3449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2781]),.i2(intermediate_reg_0[2780]),.o(intermediate_reg_1[1390])); 
fsm fsm_inst_1_3450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2779]),.i2(intermediate_reg_0[2778]),.o(intermediate_reg_1[1389])); 
mux_module mux_module_inst_1_3451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2777]),.i2(intermediate_reg_0[2776]),.o(intermediate_reg_1[1388]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2775]),.i2(intermediate_reg_0[2774]),.o(intermediate_reg_1[1387])); 
mux_module mux_module_inst_1_3453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2773]),.i2(intermediate_reg_0[2772]),.o(intermediate_reg_1[1386]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2771]),.i2(intermediate_reg_0[2770]),.o(intermediate_reg_1[1385]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2769]),.i2(intermediate_reg_0[2768]),.o(intermediate_reg_1[1384])); 
fsm fsm_inst_1_3456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2767]),.i2(intermediate_reg_0[2766]),.o(intermediate_reg_1[1383])); 
fsm fsm_inst_1_3457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2765]),.i2(intermediate_reg_0[2764]),.o(intermediate_reg_1[1382])); 
mux_module mux_module_inst_1_3458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2763]),.i2(intermediate_reg_0[2762]),.o(intermediate_reg_1[1381]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2761]),.i2(intermediate_reg_0[2760]),.o(intermediate_reg_1[1380]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2759]),.i2(intermediate_reg_0[2758]),.o(intermediate_reg_1[1379]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2757]),.i2(intermediate_reg_0[2756]),.o(intermediate_reg_1[1378]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2755]),.i2(intermediate_reg_0[2754]),.o(intermediate_reg_1[1377]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2753]),.i2(intermediate_reg_0[2752]),.o(intermediate_reg_1[1376])); 
fsm fsm_inst_1_3464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2751]),.i2(intermediate_reg_0[2750]),.o(intermediate_reg_1[1375])); 
mux_module mux_module_inst_1_3465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2749]),.i2(intermediate_reg_0[2748]),.o(intermediate_reg_1[1374]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2747]),.i2(intermediate_reg_0[2746]),.o(intermediate_reg_1[1373])); 
mux_module mux_module_inst_1_3467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2745]),.i2(intermediate_reg_0[2744]),.o(intermediate_reg_1[1372]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2743]),.i2(intermediate_reg_0[2742]),.o(intermediate_reg_1[1371])); 
fsm fsm_inst_1_3469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2741]),.i2(intermediate_reg_0[2740]),.o(intermediate_reg_1[1370])); 
mux_module mux_module_inst_1_3470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2739]),.i2(intermediate_reg_0[2738]),.o(intermediate_reg_1[1369]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2737]),.i2(intermediate_reg_0[2736]),.o(intermediate_reg_1[1368]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2735]),.i2(intermediate_reg_0[2734]),.o(intermediate_reg_1[1367]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2733]),.i2(intermediate_reg_0[2732]),.o(intermediate_reg_1[1366])); 
fsm fsm_inst_1_3474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2731]),.i2(intermediate_reg_0[2730]),.o(intermediate_reg_1[1365])); 
mux_module mux_module_inst_1_3475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2729]),.i2(intermediate_reg_0[2728]),.o(intermediate_reg_1[1364]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2727]),.i2(intermediate_reg_0[2726]),.o(intermediate_reg_1[1363])); 
mux_module mux_module_inst_1_3477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2725]),.i2(intermediate_reg_0[2724]),.o(intermediate_reg_1[1362]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2723]),.i2(intermediate_reg_0[2722]),.o(intermediate_reg_1[1361])); 
mux_module mux_module_inst_1_3479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2721]),.i2(intermediate_reg_0[2720]),.o(intermediate_reg_1[1360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2719]),.i2(intermediate_reg_0[2718]),.o(intermediate_reg_1[1359]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2717]),.i2(intermediate_reg_0[2716]),.o(intermediate_reg_1[1358])); 
mux_module mux_module_inst_1_3482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2715]),.i2(intermediate_reg_0[2714]),.o(intermediate_reg_1[1357]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2713]),.i2(intermediate_reg_0[2712]),.o(intermediate_reg_1[1356])); 
mux_module mux_module_inst_1_3484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2711]),.i2(intermediate_reg_0[2710]),.o(intermediate_reg_1[1355]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2709]),.i2(intermediate_reg_0[2708]),.o(intermediate_reg_1[1354])); 
fsm fsm_inst_1_3486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2707]),.i2(intermediate_reg_0[2706]),.o(intermediate_reg_1[1353])); 
mux_module mux_module_inst_1_3487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2705]),.i2(intermediate_reg_0[2704]),.o(intermediate_reg_1[1352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2703]),.i2(intermediate_reg_0[2702]),.o(intermediate_reg_1[1351]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2701]),.i2(intermediate_reg_0[2700]),.o(intermediate_reg_1[1350])); 
mux_module mux_module_inst_1_3490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2699]),.i2(intermediate_reg_0[2698]),.o(intermediate_reg_1[1349]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2697]),.i2(intermediate_reg_0[2696]),.o(intermediate_reg_1[1348])); 
fsm fsm_inst_1_3492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2695]),.i2(intermediate_reg_0[2694]),.o(intermediate_reg_1[1347])); 
fsm fsm_inst_1_3493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2693]),.i2(intermediate_reg_0[2692]),.o(intermediate_reg_1[1346])); 
fsm fsm_inst_1_3494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2691]),.i2(intermediate_reg_0[2690]),.o(intermediate_reg_1[1345])); 
mux_module mux_module_inst_1_3495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2689]),.i2(intermediate_reg_0[2688]),.o(intermediate_reg_1[1344]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343])); 
fsm fsm_inst_1_3497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342])); 
fsm fsm_inst_1_3498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341])); 
fsm fsm_inst_1_3499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340])); 
mux_module mux_module_inst_1_3500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338])); 
fsm fsm_inst_1_3502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337])); 
mux_module mux_module_inst_1_3503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335])); 
fsm fsm_inst_1_3505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334])); 
fsm fsm_inst_1_3506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333])); 
mux_module mux_module_inst_1_3507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330])); 
fsm fsm_inst_1_3510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329])); 
fsm fsm_inst_1_3511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328])); 
fsm fsm_inst_1_3512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327])); 
mux_module mux_module_inst_1_3513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325])); 
fsm fsm_inst_1_3515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324])); 
fsm fsm_inst_1_3516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323])); 
mux_module mux_module_inst_1_3517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321])); 
mux_module mux_module_inst_1_3519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318])); 
mux_module mux_module_inst_1_3522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316])); 
mux_module mux_module_inst_1_3524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314])); 
fsm fsm_inst_1_3526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313])); 
mux_module mux_module_inst_1_3527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310])); 
mux_module mux_module_inst_1_3530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304])); 
mux_module mux_module_inst_1_3536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301])); 
mux_module mux_module_inst_1_3539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298])); 
fsm fsm_inst_1_3542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297])); 
fsm fsm_inst_1_3543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296])); 
mux_module mux_module_inst_1_3544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291])); 
fsm fsm_inst_1_3549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290])); 
fsm fsm_inst_1_3550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289])); 
mux_module mux_module_inst_1_3551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287])); 
fsm fsm_inst_1_3553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286])); 
mux_module mux_module_inst_1_3554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284])); 
fsm fsm_inst_1_3556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283])); 
mux_module mux_module_inst_1_3557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279])); 
mux_module mux_module_inst_1_3561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275])); 
fsm fsm_inst_1_3565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274])); 
mux_module mux_module_inst_1_3566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272])); 
fsm fsm_inst_1_3568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271])); 
fsm fsm_inst_1_3569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270])); 
fsm fsm_inst_1_3570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269])); 
mux_module mux_module_inst_1_3571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267])); 
mux_module mux_module_inst_1_3573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264])); 
mux_module mux_module_inst_1_3576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262])); 
mux_module mux_module_inst_1_3578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260])); 
fsm fsm_inst_1_3580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259])); 
mux_module mux_module_inst_1_3581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257])); 
mux_module mux_module_inst_1_3583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252])); 
fsm fsm_inst_1_3588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251])); 
fsm fsm_inst_1_3589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250])); 
mux_module mux_module_inst_1_3590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247])); 
mux_module mux_module_inst_1_3593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245])); 
fsm fsm_inst_1_3595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244])); 
fsm fsm_inst_1_3596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243])); 
mux_module mux_module_inst_1_3597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241])); 
mux_module mux_module_inst_1_3599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238])); 
fsm fsm_inst_1_3602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237])); 
mux_module mux_module_inst_1_3603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234])); 
mux_module mux_module_inst_1_3606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232])); 
mux_module mux_module_inst_1_3608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230])); 
fsm fsm_inst_1_3610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229])); 
mux_module mux_module_inst_1_3611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227])); 
fsm fsm_inst_1_3613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
fsm fsm_inst_1_3614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225])); 
mux_module mux_module_inst_1_3615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222])); 
fsm fsm_inst_1_3618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221])); 
mux_module mux_module_inst_1_3619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214])); 
mux_module mux_module_inst_1_3626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212])); 
fsm fsm_inst_1_3628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211])); 
mux_module mux_module_inst_1_3629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209])); 
mux_module mux_module_inst_1_3631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206])); 
fsm fsm_inst_1_3634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205])); 
mux_module mux_module_inst_1_3635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202])); 
mux_module mux_module_inst_1_3638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198])); 
fsm fsm_inst_1_3642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197])); 
fsm fsm_inst_1_3643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196])); 
mux_module mux_module_inst_1_3644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192])); 
mux_module mux_module_inst_1_3648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190])); 
fsm fsm_inst_1_3650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189])); 
fsm fsm_inst_1_3651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188])); 
mux_module mux_module_inst_1_3652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186])); 
mux_module mux_module_inst_1_3654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180])); 
fsm fsm_inst_1_3660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179])); 
mux_module mux_module_inst_1_3661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177])); 
fsm fsm_inst_1_3663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176])); 
mux_module mux_module_inst_1_3664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174])); 
fsm fsm_inst_1_3666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173])); 
mux_module mux_module_inst_1_3667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171])); 
fsm fsm_inst_1_3669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170])); 
mux_module mux_module_inst_1_3670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167])); 
mux_module mux_module_inst_1_3673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159])); 
mux_module mux_module_inst_1_3681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
mux_module mux_module_inst_1_3683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153])); 
mux_module mux_module_inst_1_3687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150])); 
mux_module mux_module_inst_1_3690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146])); 
mux_module mux_module_inst_1_3694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144])); 
mux_module mux_module_inst_1_3696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142])); 
fsm fsm_inst_1_3698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141])); 
mux_module mux_module_inst_1_3699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136])); 
fsm fsm_inst_1_3704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135])); 
fsm fsm_inst_1_3705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134])); 
fsm fsm_inst_1_3706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133])); 
fsm fsm_inst_1_3707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132])); 
mux_module mux_module_inst_1_3708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
fsm fsm_inst_1_3710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129])); 
fsm fsm_inst_1_3711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128])); 
mux_module mux_module_inst_1_3712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
mux_module mux_module_inst_1_3715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123])); 
mux_module mux_module_inst_1_3717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121])); 
mux_module mux_module_inst_1_3719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118])); 
mux_module mux_module_inst_1_3722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115])); 
mux_module mux_module_inst_1_3725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
mux_module mux_module_inst_1_3732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106])); 
fsm fsm_inst_1_3734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
fsm fsm_inst_1_3735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
fsm fsm_inst_1_3736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
mux_module mux_module_inst_1_3737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096])); 
mux_module mux_module_inst_1_3744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094])); 
fsm fsm_inst_1_3746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
fsm fsm_inst_1_3747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
fsm fsm_inst_1_3748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
mux_module mux_module_inst_1_3749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
fsm fsm_inst_1_3751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088])); 
fsm fsm_inst_1_3752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
mux_module mux_module_inst_1_3753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
fsm fsm_inst_1_3757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082])); 
fsm fsm_inst_1_3758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081])); 
mux_module mux_module_inst_1_3759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
mux_module mux_module_inst_1_3762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076])); 
fsm fsm_inst_1_3764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075])); 
mux_module mux_module_inst_1_3765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
mux_module mux_module_inst_1_3767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069])); 
mux_module mux_module_inst_1_3771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
mux_module mux_module_inst_1_3773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065])); 
mux_module mux_module_inst_1_3775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063])); 
mux_module mux_module_inst_1_3777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058])); 
mux_module mux_module_inst_1_3782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056])); 
mux_module mux_module_inst_1_3784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
fsm fsm_inst_1_3788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051])); 
mux_module mux_module_inst_1_3789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
fsm fsm_inst_1_3793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046])); 
fsm fsm_inst_1_3794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045])); 
fsm fsm_inst_1_3795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
mux_module mux_module_inst_1_3796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
mux_module mux_module_inst_1_3798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040])); 
mux_module mux_module_inst_1_3800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
mux_module mux_module_inst_1_3809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029])); 
fsm fsm_inst_1_3811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
mux_module mux_module_inst_1_3812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
fsm fsm_inst_1_3815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024])); 
fsm fsm_inst_1_3816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
mux_module mux_module_inst_1_3817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021])); 
fsm fsm_inst_1_3819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
fsm fsm_inst_1_3820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
fsm fsm_inst_1_3821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018])); 
mux_module mux_module_inst_1_3822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
fsm fsm_inst_1_3826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013])); 
mux_module mux_module_inst_1_3827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011])); 
fsm fsm_inst_1_3829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010])); 
mux_module mux_module_inst_1_3830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008])); 
fsm fsm_inst_1_3832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
mux_module mux_module_inst_1_3833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
mux_module mux_module_inst_1_3835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
fsm fsm_inst_1_3837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
mux_module mux_module_inst_1_3838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
mux_module mux_module_inst_1_3840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
fsm fsm_inst_1_3842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
mux_module mux_module_inst_1_3843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995])); 
fsm fsm_inst_1_3845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
fsm fsm_inst_1_3846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993])); 
mux_module mux_module_inst_1_3847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
mux_module mux_module_inst_1_3852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
mux_module mux_module_inst_1_3854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
fsm fsm_inst_1_3859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
fsm fsm_inst_1_3860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
fsm fsm_inst_1_3861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978])); 
fsm fsm_inst_1_3862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
mux_module mux_module_inst_1_3863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
mux_module mux_module_inst_1_3868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
mux_module mux_module_inst_1_3871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
fsm fsm_inst_1_3873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966])); 
fsm fsm_inst_1_3874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
fsm fsm_inst_1_3875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
fsm fsm_inst_1_3876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
fsm fsm_inst_1_3877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962])); 
fsm fsm_inst_1_3878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
fsm fsm_inst_1_3879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
mux_module mux_module_inst_1_3880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
fsm fsm_inst_1_3884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
fsm fsm_inst_1_3885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954])); 
fsm fsm_inst_1_3886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
fsm fsm_inst_1_3887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
fsm fsm_inst_1_3888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
mux_module mux_module_inst_1_3889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
mux_module mux_module_inst_1_3891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947])); 
fsm fsm_inst_1_3893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
mux_module mux_module_inst_1_3894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
mux_module mux_module_inst_1_3896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
fsm fsm_inst_1_3906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
mux_module mux_module_inst_1_3907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
fsm fsm_inst_1_3909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930])); 
mux_module mux_module_inst_1_3910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
mux_module mux_module_inst_1_3913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
fsm fsm_inst_1_3915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
mux_module mux_module_inst_1_3916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
mux_module mux_module_inst_1_3922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
fsm fsm_inst_1_3927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
fsm fsm_inst_1_3928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
fsm fsm_inst_1_3929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
fsm fsm_inst_1_3930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
fsm fsm_inst_1_3931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
fsm fsm_inst_1_3932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
fsm fsm_inst_1_3933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906])); 
mux_module mux_module_inst_1_3934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
fsm fsm_inst_1_3936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
fsm fsm_inst_1_3937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
mux_module mux_module_inst_1_3938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
mux_module mux_module_inst_1_3940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
mux_module mux_module_inst_1_3942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
mux_module mux_module_inst_1_3945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
fsm fsm_inst_1_3949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
mux_module mux_module_inst_1_3950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888])); 
fsm fsm_inst_1_3952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887])); 
mux_module mux_module_inst_1_3953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
mux_module mux_module_inst_1_3957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
fsm fsm_inst_1_3959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
mux_module mux_module_inst_1_3960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
mux_module mux_module_inst_1_3964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
mux_module mux_module_inst_1_3966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
fsm fsm_inst_1_3968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
mux_module mux_module_inst_1_3969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
mux_module mux_module_inst_1_3971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
mux_module mux_module_inst_1_3973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
mux_module mux_module_inst_1_3977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
mux_module mux_module_inst_1_3979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
mux_module mux_module_inst_1_3982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
mux_module mux_module_inst_1_3984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853])); 
mux_module mux_module_inst_1_3987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851])); 
fsm fsm_inst_1_3989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
fsm fsm_inst_1_3990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
fsm fsm_inst_1_3991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
fsm fsm_inst_1_3992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
mux_module mux_module_inst_1_3993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
mux_module mux_module_inst_1_3995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
fsm fsm_inst_1_4000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
mux_module mux_module_inst_1_4001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
fsm fsm_inst_1_4003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
mux_module mux_module_inst_1_4004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
mux_module mux_module_inst_1_4007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831])); 
mux_module mux_module_inst_1_4009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
fsm fsm_inst_1_4013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
fsm fsm_inst_1_4014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
mux_module mux_module_inst_1_4015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
mux_module mux_module_inst_1_4018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
mux_module mux_module_inst_1_4020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
mux_module mux_module_inst_1_4022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
mux_module mux_module_inst_1_4024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
fsm fsm_inst_1_4026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
mux_module mux_module_inst_1_4027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
mux_module mux_module_inst_1_4029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
fsm fsm_inst_1_4031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
mux_module mux_module_inst_1_4032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
fsm fsm_inst_1_4035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
mux_module mux_module_inst_1_4036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
mux_module mux_module_inst_1_4038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
mux_module mux_module_inst_1_4040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796])); 
fsm fsm_inst_1_4044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
mux_module mux_module_inst_1_4045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
mux_module mux_module_inst_1_4048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
fsm fsm_inst_1_4051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
fsm fsm_inst_1_4052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
fsm fsm_inst_1_4053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
fsm fsm_inst_1_4054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
mux_module mux_module_inst_1_4055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
fsm fsm_inst_1_4059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
fsm fsm_inst_1_4060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
mux_module mux_module_inst_1_4061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
mux_module mux_module_inst_1_4065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
fsm fsm_inst_1_4068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
mux_module mux_module_inst_1_4069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
mux_module mux_module_inst_1_4071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
fsm fsm_inst_1_4078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
fsm fsm_inst_1_4079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
mux_module mux_module_inst_1_4080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
fsm fsm_inst_1_4082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
mux_module mux_module_inst_1_4083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
mux_module mux_module_inst_1_4086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
mux_module mux_module_inst_1_4088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
mux_module mux_module_inst_1_4090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
mux_module mux_module_inst_1_4092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
mux_module mux_module_inst_1_4100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
fsm fsm_inst_1_4103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
fsm fsm_inst_1_4104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735])); 
mux_module mux_module_inst_1_4105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
fsm fsm_inst_1_4108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
fsm fsm_inst_1_4109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
fsm fsm_inst_1_4110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729])); 
mux_module mux_module_inst_1_4111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
fsm fsm_inst_1_4114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725])); 
fsm fsm_inst_1_4115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
fsm fsm_inst_1_4116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
mux_module mux_module_inst_1_4117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
mux_module mux_module_inst_1_4120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718])); 
fsm fsm_inst_1_4122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
mux_module mux_module_inst_1_4123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
mux_module mux_module_inst_1_4125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
mux_module mux_module_inst_1_4127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
fsm fsm_inst_1_4134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
mux_module mux_module_inst_1_4135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
fsm fsm_inst_1_4137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
mux_module mux_module_inst_1_4138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
mux_module mux_module_inst_1_4140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
mux_module mux_module_inst_1_4142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
mux_module mux_module_inst_1_4144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
fsm fsm_inst_1_4149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
mux_module mux_module_inst_1_4150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
mux_module mux_module_inst_1_4152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686])); 
mux_module mux_module_inst_1_4154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
mux_module mux_module_inst_1_4157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
mux_module mux_module_inst_1_4159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
mux_module mux_module_inst_1_4161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677])); 
mux_module mux_module_inst_1_4163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
fsm fsm_inst_1_4166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
fsm fsm_inst_1_4167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
fsm fsm_inst_1_4168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671])); 
fsm fsm_inst_1_4169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
fsm fsm_inst_1_4170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
mux_module mux_module_inst_1_4171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664])); 
mux_module mux_module_inst_1_4176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
mux_module mux_module_inst_1_4178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
mux_module mux_module_inst_1_4180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
mux_module mux_module_inst_1_4182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
mux_module mux_module_inst_1_4184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653])); 
mux_module mux_module_inst_1_4187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
mux_module mux_module_inst_1_4189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
mux_module mux_module_inst_1_4191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
mux_module mux_module_inst_1_4193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
fsm fsm_inst_1_4195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
mux_module mux_module_inst_1_4196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640])); 
fsm fsm_inst_1_4200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
fsm fsm_inst_1_4201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
mux_module mux_module_inst_1_4202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635])); 
fsm fsm_inst_1_4205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
mux_module mux_module_inst_1_4206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
fsm fsm_inst_1_4210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629])); 
fsm fsm_inst_1_4211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
fsm fsm_inst_1_4212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
mux_module mux_module_inst_1_4213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
fsm fsm_inst_1_4217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
mux_module mux_module_inst_1_4218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
mux_module mux_module_inst_1_4222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
fsm fsm_inst_1_4224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
mux_module mux_module_inst_1_4225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
mux_module mux_module_inst_1_4228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
fsm fsm_inst_1_4230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
fsm fsm_inst_1_4231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
mux_module mux_module_inst_1_4232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
mux_module mux_module_inst_1_4239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599])); 
mux_module mux_module_inst_1_4241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
mux_module mux_module_inst_1_4244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_4246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
fsm fsm_inst_1_4247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
mux_module mux_module_inst_1_4248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
fsm fsm_inst_1_4251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
fsm fsm_inst_1_4252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
mux_module mux_module_inst_1_4253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
mux_module mux_module_inst_1_4260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
fsm fsm_inst_1_4263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
mux_module mux_module_inst_1_4264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
mux_module mux_module_inst_1_4267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
mux_module mux_module_inst_1_4269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
fsm fsm_inst_1_4271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
mux_module mux_module_inst_1_4272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
mux_module mux_module_inst_1_4274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
mux_module mux_module_inst_1_4278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
fsm fsm_inst_1_4280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559])); 
mux_module mux_module_inst_1_4281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_4284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
mux_module mux_module_inst_1_4285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
mux_module mux_module_inst_1_4287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
fsm fsm_inst_1_4290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
mux_module mux_module_inst_1_4291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
mux_module mux_module_inst_1_4300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
mux_module mux_module_inst_1_4302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_4305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
fsm fsm_inst_1_4306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
mux_module mux_module_inst_1_4307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531])); 
fsm fsm_inst_1_4309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530])); 
fsm fsm_inst_1_4310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
fsm fsm_inst_1_4311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
mux_module mux_module_inst_1_4312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
mux_module mux_module_inst_1_4314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523])); 
mux_module mux_module_inst_1_4317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
mux_module mux_module_inst_1_4323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
mux_module mux_module_inst_1_4326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
mux_module mux_module_inst_1_4331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
fsm fsm_inst_1_4334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
fsm fsm_inst_1_4335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
fsm fsm_inst_1_4336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
fsm fsm_inst_1_4337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
fsm fsm_inst_1_4338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
fsm fsm_inst_1_4339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
fsm fsm_inst_1_4340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
fsm fsm_inst_1_4341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
fsm fsm_inst_1_4342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
fsm fsm_inst_1_4343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
fsm fsm_inst_1_4344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
mux_module mux_module_inst_1_4345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
fsm fsm_inst_1_4347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
mux_module mux_module_inst_1_4348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
mux_module mux_module_inst_1_4359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
mux_module mux_module_inst_1_4361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_4363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
fsm fsm_inst_1_4364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
fsm fsm_inst_1_4365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
mux_module mux_module_inst_1_4366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
mux_module mux_module_inst_1_4370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462])); 
mux_module mux_module_inst_1_4378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
mux_module mux_module_inst_1_4381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
mux_module mux_module_inst_1_4383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
fsm fsm_inst_1_4388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451])); 
mux_module mux_module_inst_1_4389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
fsm fsm_inst_1_4395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
mux_module mux_module_inst_1_4396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
fsm fsm_inst_1_4399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
mux_module mux_module_inst_1_4400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
mux_module mux_module_inst_1_4405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433])); 
fsm fsm_inst_1_4407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
fsm fsm_inst_1_4408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
fsm fsm_inst_1_4409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
fsm fsm_inst_1_4410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
fsm fsm_inst_1_4411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
fsm fsm_inst_1_4412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_4413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
mux_module mux_module_inst_1_4414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
fsm fsm_inst_1_4416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
fsm fsm_inst_1_4417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
mux_module mux_module_inst_1_4418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420])); 
fsm fsm_inst_1_4420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419])); 
mux_module mux_module_inst_1_4421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
fsm fsm_inst_1_4425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
mux_module mux_module_inst_1_4426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
mux_module mux_module_inst_1_4429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
fsm fsm_inst_1_4431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
mux_module mux_module_inst_1_4432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
mux_module mux_module_inst_1_4434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404])); 
mux_module mux_module_inst_1_4436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
fsm fsm_inst_1_4438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
mux_module mux_module_inst_1_4439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
mux_module mux_module_inst_1_4441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395])); 
fsm fsm_inst_1_4445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
mux_module mux_module_inst_1_4446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392])); 
mux_module mux_module_inst_1_4448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
mux_module mux_module_inst_1_4450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387])); 
fsm fsm_inst_1_4453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386])); 
mux_module mux_module_inst_1_4454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
mux_module mux_module_inst_1_4458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
mux_module mux_module_inst_1_4461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
mux_module mux_module_inst_1_4467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
fsm fsm_inst_1_4469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370])); 
fsm fsm_inst_1_4470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
mux_module mux_module_inst_1_4471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364])); 
fsm fsm_inst_1_4476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
mux_module mux_module_inst_1_4477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361])); 
mux_module mux_module_inst_1_4479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
fsm fsm_inst_1_4483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
mux_module mux_module_inst_1_4484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351])); 
fsm fsm_inst_1_4489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
mux_module mux_module_inst_1_4490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
mux_module mux_module_inst_1_4493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
mux_module mux_module_inst_1_4496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
fsm fsm_inst_1_4498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
fsm fsm_inst_1_4499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
fsm fsm_inst_1_4500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
mux_module mux_module_inst_1_4501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
fsm fsm_inst_1_4503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
mux_module mux_module_inst_1_4504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
fsm fsm_inst_1_4506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
mux_module mux_module_inst_1_4507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
mux_module mux_module_inst_1_4512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323])); 
mux_module mux_module_inst_1_4517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
fsm fsm_inst_1_4520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
fsm fsm_inst_1_4521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318])); 
fsm fsm_inst_1_4522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317])); 
fsm fsm_inst_1_4523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316])); 
fsm fsm_inst_1_4524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
mux_module mux_module_inst_1_4525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_4529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309])); 
fsm fsm_inst_1_4531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
mux_module mux_module_inst_1_4532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
fsm fsm_inst_1_4536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
mux_module mux_module_inst_1_4537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296])); 
mux_module mux_module_inst_1_4544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
fsm fsm_inst_1_4546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
mux_module mux_module_inst_1_4547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
mux_module mux_module_inst_1_4550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
mux_module mux_module_inst_1_4552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_4559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
mux_module mux_module_inst_1_4560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
mux_module mux_module_inst_1_4563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
mux_module mux_module_inst_1_4565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
mux_module mux_module_inst_1_4567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
fsm fsm_inst_1_4570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
mux_module mux_module_inst_1_4571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
fsm fsm_inst_1_4574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
fsm fsm_inst_1_4575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
mux_module mux_module_inst_1_4576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
fsm fsm_inst_1_4581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
mux_module mux_module_inst_1_4582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
fsm fsm_inst_1_4585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
fsm fsm_inst_1_4586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
mux_module mux_module_inst_1_4587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
fsm fsm_inst_1_4589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
mux_module mux_module_inst_1_4590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247])); 
fsm fsm_inst_1_4593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
mux_module mux_module_inst_1_4594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
fsm fsm_inst_1_4597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
fsm fsm_inst_1_4598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241])); 
mux_module mux_module_inst_1_4599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
mux_module mux_module_inst_1_4602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
fsm fsm_inst_1_4605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
mux_module mux_module_inst_1_4606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
fsm fsm_inst_1_4608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
fsm fsm_inst_1_4609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
mux_module mux_module_inst_1_4610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
fsm fsm_inst_1_4612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
fsm fsm_inst_1_4613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
fsm fsm_inst_1_4614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
fsm fsm_inst_1_4615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
fsm fsm_inst_1_4616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
fsm fsm_inst_1_4617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
mux_module mux_module_inst_1_4618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
mux_module mux_module_inst_1_4620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
mux_module mux_module_inst_1_4622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
fsm fsm_inst_1_4625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
fsm fsm_inst_1_4626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
mux_module mux_module_inst_1_4627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
mux_module mux_module_inst_1_4630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
mux_module mux_module_inst_1_4633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
mux_module mux_module_inst_1_4635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
fsm fsm_inst_1_4638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
mux_module mux_module_inst_1_4639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
fsm fsm_inst_1_4641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_4642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
mux_module mux_module_inst_1_4645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
fsm fsm_inst_1_4647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
mux_module mux_module_inst_1_4648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
fsm fsm_inst_1_4650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
mux_module mux_module_inst_1_4651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
fsm fsm_inst_1_4653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
fsm fsm_inst_1_4654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185])); 
fsm fsm_inst_1_4655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
mux_module mux_module_inst_1_4656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
mux_module mux_module_inst_1_4658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
fsm fsm_inst_1_4660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
mux_module mux_module_inst_1_4661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177])); 
mux_module mux_module_inst_1_4663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
fsm fsm_inst_1_4665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
fsm fsm_inst_1_4666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
fsm fsm_inst_1_4667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
fsm fsm_inst_1_4668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
mux_module mux_module_inst_1_4669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
fsm fsm_inst_1_4672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167])); 
mux_module mux_module_inst_1_4673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
fsm fsm_inst_1_4675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
fsm fsm_inst_1_4676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
mux_module mux_module_inst_1_4677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
fsm fsm_inst_1_4680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
fsm fsm_inst_1_4681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
mux_module mux_module_inst_1_4682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
fsm fsm_inst_1_4684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
fsm fsm_inst_1_4685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
mux_module mux_module_inst_1_4686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
fsm fsm_inst_1_4689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
mux_module mux_module_inst_1_4690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
mux_module mux_module_inst_1_4692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
fsm fsm_inst_1_4694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
mux_module mux_module_inst_1_4695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
fsm fsm_inst_1_4697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_4698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
mux_module mux_module_inst_1_4699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
mux_module mux_module_inst_1_4701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
fsm fsm_inst_1_4703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
fsm fsm_inst_1_4704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
mux_module mux_module_inst_1_4705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
mux_module mux_module_inst_1_4707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
mux_module mux_module_inst_1_4711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
mux_module mux_module_inst_1_4714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123])); 
mux_module mux_module_inst_1_4717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
mux_module mux_module_inst_1_4721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
mux_module mux_module_inst_1_4724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
fsm fsm_inst_1_4726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
mux_module mux_module_inst_1_4727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
fsm fsm_inst_1_4730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
mux_module mux_module_inst_1_4731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
fsm fsm_inst_1_4733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
mux_module mux_module_inst_1_4734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
mux_module mux_module_inst_1_4736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
mux_module mux_module_inst_1_4741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
mux_module mux_module_inst_1_4744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
fsm fsm_inst_1_4748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
fsm fsm_inst_1_4749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
mux_module mux_module_inst_1_4750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
mux_module mux_module_inst_1_4752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
mux_module mux_module_inst_1_4754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
mux_module mux_module_inst_1_4759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77])); 
fsm fsm_inst_1_4763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
mux_module mux_module_inst_1_4764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
fsm fsm_inst_1_4769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
mux_module mux_module_inst_1_4770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_4774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
mux_module mux_module_inst_1_4780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
fsm fsm_inst_1_4782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57])); 
fsm fsm_inst_1_4783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
fsm fsm_inst_1_4784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
fsm fsm_inst_1_4785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
mux_module mux_module_inst_1_4786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52])); 
fsm fsm_inst_1_4788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
fsm fsm_inst_1_4789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_4790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
mux_module mux_module_inst_1_4791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
fsm fsm_inst_1_4794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
fsm fsm_inst_1_4795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
fsm fsm_inst_1_4796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
fsm fsm_inst_1_4797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
fsm fsm_inst_1_4798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_4799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38])); 
fsm fsm_inst_1_4802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
mux_module mux_module_inst_1_4803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
mux_module mux_module_inst_1_4809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
fsm fsm_inst_1_4815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
mux_module mux_module_inst_1_4816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
fsm fsm_inst_1_4820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
fsm fsm_inst_1_4821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18])); 
fsm fsm_inst_1_4822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
mux_module mux_module_inst_1_4823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_4825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
fsm fsm_inst_1_4828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
fsm fsm_inst_1_4829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
fsm fsm_inst_1_4830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9])); 
mux_module mux_module_inst_1_4831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
fsm fsm_inst_1_4833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
mux_module mux_module_inst_1_4834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
fsm fsm_inst_1_4836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
fsm fsm_inst_1_4837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
fsm fsm_inst_1_4838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
mux_module mux_module_inst_1_4839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
always@(posedge clk) begin 
outp [4839:0] <= intermediate_reg_1; 
outp[9599:4840] <= intermediate_reg_1[4759:0] ; 
end 
endmodule 
 

module interface_24(input reg [4319:0] inp, output reg [5119:0] outp, input clk, input reset);
always@(posedge clk) begin 
outp[4319:0] <= inp ; 
outp[5119:4320] <= inp[799:0] ; 
end 
endmodule 

module interface_25(input reg [2239:0] inp, output reg [527:0] outp, input clk, input reset);
reg [2239:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1119:0]intermediate_reg_1; 
 
fsm fsm_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111])); 
mux_module mux_module_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
mux_module mux_module_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
fsm fsm_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094])); 
fsm fsm_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
fsm fsm_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086])); 
fsm fsm_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084])); 
fsm fsm_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
mux_module mux_module_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071])); 
mux_module mux_module_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069])); 
fsm fsm_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068])); 
fsm fsm_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
fsm fsm_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066])); 
fsm fsm_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059])); 
fsm fsm_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058])); 
fsm fsm_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057])); 
mux_module mux_module_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055])); 
fsm fsm_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
mux_module mux_module_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046])); 
fsm fsm_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045])); 
fsm fsm_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044])); 
fsm fsm_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041])); 
mux_module mux_module_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032])); 
fsm fsm_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
mux_module mux_module_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027])); 
fsm fsm_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026])); 
fsm fsm_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016])); 
fsm fsm_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014])); 
mux_module mux_module_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003])); 
fsm fsm_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001])); 
fsm fsm_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991])); 
fsm fsm_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990])); 
fsm fsm_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
mux_module mux_module_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
fsm fsm_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
fsm fsm_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
fsm fsm_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978])); 
fsm fsm_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
fsm fsm_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
fsm fsm_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
mux_module mux_module_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962])); 
fsm fsm_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
mux_module mux_module_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
mux_module mux_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950])); 
mux_module mux_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
mux_module mux_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
fsm fsm_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940])); 
fsm fsm_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
fsm fsm_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925])); 
fsm fsm_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
mux_module mux_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
mux_module mux_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911])); 
mux_module mux_module_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
fsm fsm_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
mux_module mux_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906])); 
fsm fsm_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
fsm fsm_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
fsm fsm_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
fsm fsm_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891])); 
fsm fsm_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
fsm fsm_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
mux_module mux_module_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
fsm fsm_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
fsm fsm_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
mux_module mux_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
mux_module mux_module_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876])); 
fsm fsm_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
fsm fsm_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873])); 
fsm fsm_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
fsm fsm_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
fsm fsm_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
mux_module mux_module_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
mux_module mux_module_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
fsm fsm_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829])); 
fsm fsm_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
fsm fsm_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
mux_module mux_module_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
mux_module mux_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
fsm fsm_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
fsm fsm_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
fsm fsm_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815])); 
fsm fsm_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
fsm fsm_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
fsm fsm_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800])); 
fsm fsm_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
fsm fsm_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
fsm fsm_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
fsm fsm_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
fsm fsm_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
fsm fsm_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
fsm fsm_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773])); 
mux_module mux_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
fsm fsm_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770])); 
fsm fsm_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
fsm fsm_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
mux_module mux_module_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761])); 
fsm fsm_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
fsm fsm_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
fsm fsm_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757])); 
mux_module mux_module_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755])); 
fsm fsm_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754])); 
fsm fsm_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753])); 
mux_module mux_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
fsm fsm_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
mux_module mux_module_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
fsm fsm_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
mux_module mux_module_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
fsm fsm_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
fsm fsm_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
mux_module mux_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733])); 
fsm fsm_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732])); 
mux_module mux_module_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
fsm fsm_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
fsm fsm_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
fsm fsm_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
mux_module mux_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
fsm fsm_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
fsm fsm_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
fsm fsm_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
fsm fsm_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
mux_module mux_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
mux_module mux_module_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700])); 
fsm fsm_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
fsm fsm_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698])); 
fsm fsm_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697])); 
mux_module mux_module_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
mux_module mux_module_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
fsm fsm_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
fsm fsm_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
fsm fsm_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
fsm fsm_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687])); 
mux_module mux_module_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683])); 
fsm fsm_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682])); 
fsm fsm_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
fsm fsm_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
mux_module mux_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
fsm fsm_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
fsm fsm_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
mux_module mux_module_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
fsm fsm_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
mux_module mux_module_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654])); 
mux_module mux_module_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
fsm fsm_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
mux_module mux_module_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
fsm fsm_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
mux_module mux_module_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
mux_module mux_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
fsm fsm_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633])); 
fsm fsm_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632])); 
fsm fsm_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
fsm fsm_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
fsm fsm_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
mux_module mux_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
fsm fsm_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
mux_module mux_module_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
fsm fsm_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
mux_module mux_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
fsm fsm_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
fsm fsm_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
mux_module mux_module_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
mux_module mux_module_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
fsm fsm_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
fsm fsm_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567])); 
mux_module mux_module_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
fsm fsm_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
fsm fsm_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
mux_module mux_module_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
fsm fsm_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
mux_module mux_module_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
mux_module mux_module_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528])); 
mux_module mux_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516])); 
mux_module mux_module_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503])); 
fsm fsm_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
fsm fsm_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
mux_module mux_module_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
fsm fsm_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
mux_module mux_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487])); 
fsm fsm_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
mux_module mux_module_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
fsm fsm_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
mux_module mux_module_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
fsm fsm_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474])); 
fsm fsm_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
fsm fsm_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469])); 
fsm fsm_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
fsm fsm_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457])); 
fsm fsm_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
fsm fsm_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
mux_module mux_module_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
fsm fsm_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447])); 
mux_module mux_module_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
fsm fsm_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
mux_module mux_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
fsm fsm_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430])); 
fsm fsm_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
mux_module mux_module_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425])); 
mux_module mux_module_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
mux_module mux_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
mux_module mux_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
fsm fsm_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
mux_module mux_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
fsm fsm_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
fsm fsm_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373])); 
fsm fsm_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
mux_module mux_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
fsm fsm_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
fsm fsm_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
mux_module mux_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
fsm fsm_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349])); 
fsm fsm_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
fsm fsm_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347])); 
fsm fsm_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
fsm fsm_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
mux_module mux_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
fsm fsm_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342])); 
fsm fsm_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
mux_module mux_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337])); 
fsm fsm_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
mux_module mux_module_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
mux_module mux_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
mux_module mux_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
mux_module mux_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
fsm fsm_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
fsm fsm_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314])); 
fsm fsm_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
fsm fsm_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
fsm fsm_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308])); 
fsm fsm_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
fsm fsm_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
mux_module mux_module_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
mux_module mux_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
fsm fsm_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297])); 
mux_module mux_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295])); 
fsm fsm_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
fsm fsm_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
fsm fsm_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
mux_module mux_module_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
fsm fsm_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
fsm fsm_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
fsm fsm_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
mux_module mux_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
fsm fsm_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
mux_module mux_module_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
mux_module mux_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
mux_module mux_module_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
mux_module mux_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
mux_module mux_module_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
fsm fsm_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
mux_module mux_module_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
mux_module mux_module_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
mux_module mux_module_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255])); 
fsm fsm_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254])); 
mux_module mux_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
mux_module mux_module_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
mux_module mux_module_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246])); 
fsm fsm_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
fsm fsm_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
fsm fsm_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
fsm fsm_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
fsm fsm_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
fsm fsm_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
mux_module mux_module_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
mux_module mux_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
fsm fsm_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
fsm fsm_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
mux_module mux_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
mux_module mux_module_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
mux_module mux_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
fsm fsm_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219])); 
fsm fsm_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
fsm fsm_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
fsm fsm_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
fsm fsm_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
fsm fsm_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
mux_module mux_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
mux_module mux_module_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
mux_module mux_module_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
fsm fsm_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195])); 
fsm fsm_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
mux_module mux_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
mux_module mux_module_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
mux_module mux_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
mux_module mux_module_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181])); 
fsm fsm_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180])); 
fsm fsm_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
fsm fsm_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
mux_module mux_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
fsm fsm_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
mux_module mux_module_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
mux_module mux_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
mux_module mux_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
mux_module mux_module_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
mux_module mux_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
fsm fsm_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
fsm fsm_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158])); 
fsm fsm_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
mux_module mux_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155])); 
mux_module mux_module_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152])); 
fsm fsm_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
fsm fsm_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
mux_module mux_module_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
fsm fsm_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
mux_module mux_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
fsm fsm_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
fsm fsm_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137])); 
fsm fsm_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
mux_module mux_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
fsm fsm_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
mux_module mux_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
fsm fsm_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
mux_module mux_module_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
fsm fsm_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
fsm fsm_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
mux_module mux_module_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121])); 
mux_module mux_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
mux_module mux_module_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
fsm fsm_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
mux_module mux_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
fsm fsm_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
fsm fsm_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
fsm fsm_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108])); 
mux_module mux_module_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
fsm fsm_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104])); 
fsm fsm_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
fsm fsm_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
fsm fsm_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95])); 
fsm fsm_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
fsm fsm_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93])); 
mux_module mux_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88])); 
fsm fsm_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87])); 
mux_module mux_module_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
mux_module mux_module_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
mux_module mux_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
mux_module mux_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
mux_module mux_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
fsm fsm_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71])); 
mux_module mux_module_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
fsm fsm_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68])); 
mux_module mux_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64])); 
mux_module mux_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62])); 
fsm fsm_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
fsm fsm_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
fsm fsm_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
mux_module mux_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56])); 
mux_module mux_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54])); 
mux_module mux_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
mux_module mux_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
mux_module mux_module_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
mux_module mux_module_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
mux_module mux_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37])); 
fsm fsm_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36])); 
fsm fsm_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
fsm fsm_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
mux_module mux_module_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
fsm fsm_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
fsm fsm_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
fsm fsm_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
fsm fsm_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
mux_module mux_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
mux_module mux_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
fsm fsm_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
fsm fsm_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13])); 
mux_module mux_module_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
mux_module mux_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
fsm fsm_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
fsm fsm_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
fsm fsm_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
mux_module mux_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
reg [559:0]intermediate_reg_2; 
 
fsm fsm_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1119]),.i2(intermediate_reg_1[1118]),.o(intermediate_reg_2[559])); 
mux_module mux_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1117]),.i2(intermediate_reg_1[1116]),.o(intermediate_reg_2[558]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1115]),.i2(intermediate_reg_1[1114]),.o(intermediate_reg_2[557])); 
fsm fsm_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1113]),.i2(intermediate_reg_1[1112]),.o(intermediate_reg_2[556])); 
mux_module mux_module_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1111]),.i2(intermediate_reg_1[1110]),.o(intermediate_reg_2[555]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1109]),.i2(intermediate_reg_1[1108]),.o(intermediate_reg_2[554]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1107]),.i2(intermediate_reg_1[1106]),.o(intermediate_reg_2[553])); 
fsm fsm_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1105]),.i2(intermediate_reg_1[1104]),.o(intermediate_reg_2[552])); 
mux_module mux_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1103]),.i2(intermediate_reg_1[1102]),.o(intermediate_reg_2[551]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1101]),.i2(intermediate_reg_1[1100]),.o(intermediate_reg_2[550]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1099]),.i2(intermediate_reg_1[1098]),.o(intermediate_reg_2[549]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1097]),.i2(intermediate_reg_1[1096]),.o(intermediate_reg_2[548]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1095]),.i2(intermediate_reg_1[1094]),.o(intermediate_reg_2[547]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1093]),.i2(intermediate_reg_1[1092]),.o(intermediate_reg_2[546])); 
mux_module mux_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1091]),.i2(intermediate_reg_1[1090]),.o(intermediate_reg_2[545]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1089]),.i2(intermediate_reg_1[1088]),.o(intermediate_reg_2[544])); 
mux_module mux_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1087]),.i2(intermediate_reg_1[1086]),.o(intermediate_reg_2[543]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1085]),.i2(intermediate_reg_1[1084]),.o(intermediate_reg_2[542]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1083]),.i2(intermediate_reg_1[1082]),.o(intermediate_reg_2[541]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1081]),.i2(intermediate_reg_1[1080]),.o(intermediate_reg_2[540])); 
fsm fsm_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1079]),.i2(intermediate_reg_1[1078]),.o(intermediate_reg_2[539])); 
fsm fsm_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1077]),.i2(intermediate_reg_1[1076]),.o(intermediate_reg_2[538])); 
fsm fsm_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1075]),.i2(intermediate_reg_1[1074]),.o(intermediate_reg_2[537])); 
mux_module mux_module_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1073]),.i2(intermediate_reg_1[1072]),.o(intermediate_reg_2[536]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1071]),.i2(intermediate_reg_1[1070]),.o(intermediate_reg_2[535])); 
mux_module mux_module_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1069]),.i2(intermediate_reg_1[1068]),.o(intermediate_reg_2[534]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1067]),.i2(intermediate_reg_1[1066]),.o(intermediate_reg_2[533])); 
fsm fsm_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1065]),.i2(intermediate_reg_1[1064]),.o(intermediate_reg_2[532])); 
mux_module mux_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1063]),.i2(intermediate_reg_1[1062]),.o(intermediate_reg_2[531]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1061]),.i2(intermediate_reg_1[1060]),.o(intermediate_reg_2[530])); 
fsm fsm_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1059]),.i2(intermediate_reg_1[1058]),.o(intermediate_reg_2[529])); 
fsm fsm_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1057]),.i2(intermediate_reg_1[1056]),.o(intermediate_reg_2[528])); 
mux_module mux_module_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1055]),.i2(intermediate_reg_1[1054]),.o(intermediate_reg_2[527]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1053]),.i2(intermediate_reg_1[1052]),.o(intermediate_reg_2[526])); 
mux_module mux_module_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1051]),.i2(intermediate_reg_1[1050]),.o(intermediate_reg_2[525]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1049]),.i2(intermediate_reg_1[1048]),.o(intermediate_reg_2[524])); 
mux_module mux_module_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1047]),.i2(intermediate_reg_1[1046]),.o(intermediate_reg_2[523]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1045]),.i2(intermediate_reg_1[1044]),.o(intermediate_reg_2[522]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1043]),.i2(intermediate_reg_1[1042]),.o(intermediate_reg_2[521]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1041]),.i2(intermediate_reg_1[1040]),.o(intermediate_reg_2[520])); 
mux_module mux_module_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1039]),.i2(intermediate_reg_1[1038]),.o(intermediate_reg_2[519]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1037]),.i2(intermediate_reg_1[1036]),.o(intermediate_reg_2[518]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1035]),.i2(intermediate_reg_1[1034]),.o(intermediate_reg_2[517])); 
fsm fsm_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1033]),.i2(intermediate_reg_1[1032]),.o(intermediate_reg_2[516])); 
mux_module mux_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1031]),.i2(intermediate_reg_1[1030]),.o(intermediate_reg_2[515]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1029]),.i2(intermediate_reg_1[1028]),.o(intermediate_reg_2[514]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513])); 
fsm fsm_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512])); 
fsm fsm_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511])); 
fsm fsm_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510])); 
mux_module mux_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508])); 
mux_module mux_module_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506])); 
mux_module mux_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502])); 
mux_module mux_module_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500])); 
mux_module mux_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498])); 
mux_module mux_module_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495])); 
fsm fsm_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494])); 
fsm fsm_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493])); 
fsm fsm_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492])); 
fsm fsm_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491])); 
fsm fsm_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490])); 
mux_module mux_module_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487])); 
mux_module mux_module_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485])); 
fsm fsm_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484])); 
mux_module mux_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482])); 
fsm fsm_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481])); 
mux_module mux_module_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
mux_module mux_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475])); 
mux_module mux_module_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473])); 
fsm fsm_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472])); 
fsm fsm_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471])); 
fsm fsm_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470])); 
mux_module mux_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467])); 
fsm fsm_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466])); 
mux_module mux_module_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461])); 
mux_module mux_module_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459])); 
fsm fsm_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458])); 
mux_module mux_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453])); 
mux_module mux_module_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450])); 
fsm fsm_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449])); 
fsm fsm_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448])); 
fsm fsm_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447])); 
mux_module mux_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443])); 
fsm fsm_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442])); 
fsm fsm_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441])); 
mux_module mux_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437])); 
fsm fsm_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436])); 
fsm fsm_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435])); 
mux_module mux_module_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433])); 
mux_module mux_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431])); 
mux_module mux_module_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428])); 
mux_module mux_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420])); 
fsm fsm_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419])); 
fsm fsm_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418])); 
mux_module mux_module_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415])); 
fsm fsm_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414])); 
mux_module mux_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412])); 
fsm fsm_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411])); 
mux_module mux_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408])); 
fsm fsm_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407])); 
fsm fsm_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406])); 
fsm fsm_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405])); 
fsm fsm_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404])); 
fsm fsm_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403])); 
mux_module mux_module_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401])); 
mux_module mux_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399])); 
mux_module mux_module_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397])); 
mux_module mux_module_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393])); 
fsm fsm_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392])); 
fsm fsm_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391])); 
fsm fsm_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390])); 
fsm fsm_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389])); 
mux_module mux_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384])); 
mux_module mux_module_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382])); 
fsm fsm_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
fsm fsm_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
fsm fsm_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379])); 
fsm fsm_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378])); 
fsm fsm_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377])); 
mux_module mux_module_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375])); 
mux_module mux_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373])); 
mux_module mux_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370])); 
mux_module mux_module_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367])); 
mux_module mux_module_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365])); 
fsm fsm_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364])); 
fsm fsm_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363])); 
fsm fsm_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362])); 
fsm fsm_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361])); 
fsm fsm_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360])); 
fsm fsm_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359])); 
fsm fsm_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
mux_module mux_module_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354])); 
mux_module mux_module_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351])); 
fsm fsm_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350])); 
fsm fsm_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349])); 
fsm fsm_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348])); 
fsm fsm_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
mux_module mux_module_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345])); 
fsm fsm_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
mux_module mux_module_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342])); 
mux_module mux_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336])); 
fsm fsm_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
fsm fsm_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334])); 
fsm fsm_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333])); 
fsm fsm_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332])); 
fsm fsm_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331])); 
fsm fsm_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330])); 
fsm fsm_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
mux_module mux_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327])); 
fsm fsm_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326])); 
mux_module mux_module_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324])); 
fsm fsm_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323])); 
fsm fsm_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322])); 
fsm fsm_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321])); 
fsm fsm_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320])); 
mux_module mux_module_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318])); 
fsm fsm_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317])); 
mux_module mux_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315])); 
fsm fsm_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314])); 
mux_module mux_module_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310])); 
mux_module mux_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307])); 
mux_module mux_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305])); 
mux_module mux_module_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302])); 
fsm fsm_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
mux_module mux_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297])); 
mux_module mux_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
mux_module mux_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
mux_module mux_module_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289])); 
mux_module mux_module_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287])); 
fsm fsm_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286])); 
fsm fsm_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285])); 
mux_module mux_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283])); 
mux_module mux_module_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276])); 
mux_module mux_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274])); 
fsm fsm_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
mux_module mux_module_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
fsm fsm_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270])); 
mux_module mux_module_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268])); 
mux_module mux_module_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265])); 
mux_module mux_module_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
fsm fsm_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261])); 
fsm fsm_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
mux_module mux_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257])); 
mux_module mux_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255])); 
mux_module mux_module_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252])); 
mux_module mux_module_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
mux_module mux_module_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247])); 
mux_module mux_module_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
fsm fsm_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244])); 
fsm fsm_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243])); 
mux_module mux_module_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241])); 
fsm fsm_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240])); 
mux_module mux_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
fsm fsm_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
mux_module mux_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231])); 
fsm fsm_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230])); 
mux_module mux_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
mux_module mux_module_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
mux_module mux_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223])); 
mux_module mux_module_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218])); 
mux_module mux_module_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
mux_module mux_module_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
fsm fsm_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210])); 
fsm fsm_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209])); 
fsm fsm_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208])); 
fsm fsm_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
mux_module mux_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204])); 
fsm fsm_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203])); 
mux_module mux_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197])); 
fsm fsm_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
fsm fsm_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195])); 
fsm fsm_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194])); 
mux_module mux_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192])); 
fsm fsm_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191])); 
fsm fsm_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190])); 
mux_module mux_module_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
fsm fsm_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187])); 
mux_module mux_module_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184])); 
mux_module mux_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180])); 
fsm fsm_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179])); 
fsm fsm_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178])); 
fsm fsm_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177])); 
fsm fsm_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176])); 
mux_module mux_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
fsm fsm_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172])); 
fsm fsm_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
mux_module mux_module_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169])); 
fsm fsm_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168])); 
fsm fsm_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167])); 
mux_module mux_module_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165])); 
fsm fsm_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164])); 
fsm fsm_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
mux_module mux_module_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160])); 
fsm fsm_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
fsm fsm_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158])); 
mux_module mux_module_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156])); 
fsm fsm_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155])); 
fsm fsm_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154])); 
fsm fsm_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153])); 
mux_module mux_module_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
mux_module mux_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148])); 
fsm fsm_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147])); 
mux_module mux_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145])); 
fsm fsm_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144])); 
mux_module mux_module_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141])); 
mux_module mux_module_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
mux_module mux_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
fsm fsm_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133])); 
mux_module mux_module_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131])); 
mux_module mux_module_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
fsm fsm_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126])); 
fsm fsm_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
fsm fsm_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124])); 
mux_module mux_module_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120])); 
mux_module mux_module_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118])); 
mux_module mux_module_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
fsm fsm_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113])); 
mux_module mux_module_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110])); 
fsm fsm_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
mux_module mux_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103])); 
fsm fsm_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102])); 
mux_module mux_module_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99])); 
mux_module mux_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
mux_module mux_module_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94])); 
fsm fsm_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
mux_module mux_module_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
mux_module mux_module_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88])); 
fsm fsm_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
mux_module mux_module_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85])); 
fsm fsm_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
mux_module mux_module_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82])); 
mux_module mux_module_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80])); 
mux_module mux_module_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
mux_module mux_module_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72])); 
mux_module mux_module_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70])); 
mux_module mux_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66])); 
mux_module mux_module_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62])); 
fsm fsm_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
mux_module mux_module_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58])); 
mux_module mux_module_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56])); 
fsm fsm_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55])); 
mux_module mux_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
mux_module mux_module_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50])); 
mux_module mux_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48])); 
mux_module mux_module_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44])); 
fsm fsm_inst_2_516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
fsm fsm_inst_2_517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42])); 
mux_module mux_module_inst_2_518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
mux_module mux_module_inst_2_523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34])); 
mux_module mux_module_inst_2_526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31])); 
mux_module mux_module_inst_2_529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29])); 
fsm fsm_inst_2_531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
fsm fsm_inst_2_532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27])); 
fsm fsm_inst_2_533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26])); 
mux_module mux_module_inst_2_534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23])); 
mux_module mux_module_inst_2_537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17])); 
mux_module mux_module_inst_2_543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15])); 
fsm fsm_inst_2_545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14])); 
mux_module mux_module_inst_2_546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11])); 
fsm fsm_inst_2_549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10])); 
mux_module mux_module_inst_2_550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8])); 
fsm fsm_inst_2_552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
fsm fsm_inst_2_553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6])); 
mux_module mux_module_inst_2_554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2])); 
fsm fsm_inst_2_558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
mux_module mux_module_inst_2_559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0]),.sel(intermediate_reg_1[0])); 
reg [279:0]intermediate_reg_3; 
 
mux_module mux_module_inst_3_0(.clk(clk),.reset(reset),.i1(intermediate_reg_2[559]),.i2(intermediate_reg_2[558]),.o(intermediate_reg_3[279]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_1(.clk(clk),.reset(reset),.i1(intermediate_reg_2[557]),.i2(intermediate_reg_2[556]),.o(intermediate_reg_3[278])); 
mux_module mux_module_inst_3_2(.clk(clk),.reset(reset),.i1(intermediate_reg_2[555]),.i2(intermediate_reg_2[554]),.o(intermediate_reg_3[277]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_3(.clk(clk),.reset(reset),.i1(intermediate_reg_2[553]),.i2(intermediate_reg_2[552]),.o(intermediate_reg_3[276])); 
fsm fsm_inst_3_4(.clk(clk),.reset(reset),.i1(intermediate_reg_2[551]),.i2(intermediate_reg_2[550]),.o(intermediate_reg_3[275])); 
mux_module mux_module_inst_3_5(.clk(clk),.reset(reset),.i1(intermediate_reg_2[549]),.i2(intermediate_reg_2[548]),.o(intermediate_reg_3[274]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_6(.clk(clk),.reset(reset),.i1(intermediate_reg_2[547]),.i2(intermediate_reg_2[546]),.o(intermediate_reg_3[273]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_7(.clk(clk),.reset(reset),.i1(intermediate_reg_2[545]),.i2(intermediate_reg_2[544]),.o(intermediate_reg_3[272])); 
fsm fsm_inst_3_8(.clk(clk),.reset(reset),.i1(intermediate_reg_2[543]),.i2(intermediate_reg_2[542]),.o(intermediate_reg_3[271])); 
mux_module mux_module_inst_3_9(.clk(clk),.reset(reset),.i1(intermediate_reg_2[541]),.i2(intermediate_reg_2[540]),.o(intermediate_reg_3[270]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_10(.clk(clk),.reset(reset),.i1(intermediate_reg_2[539]),.i2(intermediate_reg_2[538]),.o(intermediate_reg_3[269]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_11(.clk(clk),.reset(reset),.i1(intermediate_reg_2[537]),.i2(intermediate_reg_2[536]),.o(intermediate_reg_3[268])); 
mux_module mux_module_inst_3_12(.clk(clk),.reset(reset),.i1(intermediate_reg_2[535]),.i2(intermediate_reg_2[534]),.o(intermediate_reg_3[267]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_13(.clk(clk),.reset(reset),.i1(intermediate_reg_2[533]),.i2(intermediate_reg_2[532]),.o(intermediate_reg_3[266])); 
mux_module mux_module_inst_3_14(.clk(clk),.reset(reset),.i1(intermediate_reg_2[531]),.i2(intermediate_reg_2[530]),.o(intermediate_reg_3[265]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_15(.clk(clk),.reset(reset),.i1(intermediate_reg_2[529]),.i2(intermediate_reg_2[528]),.o(intermediate_reg_3[264]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_16(.clk(clk),.reset(reset),.i1(intermediate_reg_2[527]),.i2(intermediate_reg_2[526]),.o(intermediate_reg_3[263])); 
mux_module mux_module_inst_3_17(.clk(clk),.reset(reset),.i1(intermediate_reg_2[525]),.i2(intermediate_reg_2[524]),.o(intermediate_reg_3[262]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_18(.clk(clk),.reset(reset),.i1(intermediate_reg_2[523]),.i2(intermediate_reg_2[522]),.o(intermediate_reg_3[261]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_19(.clk(clk),.reset(reset),.i1(intermediate_reg_2[521]),.i2(intermediate_reg_2[520]),.o(intermediate_reg_3[260]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_20(.clk(clk),.reset(reset),.i1(intermediate_reg_2[519]),.i2(intermediate_reg_2[518]),.o(intermediate_reg_3[259]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_21(.clk(clk),.reset(reset),.i1(intermediate_reg_2[517]),.i2(intermediate_reg_2[516]),.o(intermediate_reg_3[258]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_22(.clk(clk),.reset(reset),.i1(intermediate_reg_2[515]),.i2(intermediate_reg_2[514]),.o(intermediate_reg_3[257])); 
mux_module mux_module_inst_3_23(.clk(clk),.reset(reset),.i1(intermediate_reg_2[513]),.i2(intermediate_reg_2[512]),.o(intermediate_reg_3[256]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_24(.clk(clk),.reset(reset),.i1(intermediate_reg_2[511]),.i2(intermediate_reg_2[510]),.o(intermediate_reg_3[255]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_25(.clk(clk),.reset(reset),.i1(intermediate_reg_2[509]),.i2(intermediate_reg_2[508]),.o(intermediate_reg_3[254]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_26(.clk(clk),.reset(reset),.i1(intermediate_reg_2[507]),.i2(intermediate_reg_2[506]),.o(intermediate_reg_3[253]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_27(.clk(clk),.reset(reset),.i1(intermediate_reg_2[505]),.i2(intermediate_reg_2[504]),.o(intermediate_reg_3[252]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_28(.clk(clk),.reset(reset),.i1(intermediate_reg_2[503]),.i2(intermediate_reg_2[502]),.o(intermediate_reg_3[251]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_29(.clk(clk),.reset(reset),.i1(intermediate_reg_2[501]),.i2(intermediate_reg_2[500]),.o(intermediate_reg_3[250])); 
mux_module mux_module_inst_3_30(.clk(clk),.reset(reset),.i1(intermediate_reg_2[499]),.i2(intermediate_reg_2[498]),.o(intermediate_reg_3[249]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_31(.clk(clk),.reset(reset),.i1(intermediate_reg_2[497]),.i2(intermediate_reg_2[496]),.o(intermediate_reg_3[248]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_32(.clk(clk),.reset(reset),.i1(intermediate_reg_2[495]),.i2(intermediate_reg_2[494]),.o(intermediate_reg_3[247])); 
mux_module mux_module_inst_3_33(.clk(clk),.reset(reset),.i1(intermediate_reg_2[493]),.i2(intermediate_reg_2[492]),.o(intermediate_reg_3[246]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_34(.clk(clk),.reset(reset),.i1(intermediate_reg_2[491]),.i2(intermediate_reg_2[490]),.o(intermediate_reg_3[245]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_35(.clk(clk),.reset(reset),.i1(intermediate_reg_2[489]),.i2(intermediate_reg_2[488]),.o(intermediate_reg_3[244])); 
fsm fsm_inst_3_36(.clk(clk),.reset(reset),.i1(intermediate_reg_2[487]),.i2(intermediate_reg_2[486]),.o(intermediate_reg_3[243])); 
fsm fsm_inst_3_37(.clk(clk),.reset(reset),.i1(intermediate_reg_2[485]),.i2(intermediate_reg_2[484]),.o(intermediate_reg_3[242])); 
mux_module mux_module_inst_3_38(.clk(clk),.reset(reset),.i1(intermediate_reg_2[483]),.i2(intermediate_reg_2[482]),.o(intermediate_reg_3[241]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_39(.clk(clk),.reset(reset),.i1(intermediate_reg_2[481]),.i2(intermediate_reg_2[480]),.o(intermediate_reg_3[240])); 
mux_module mux_module_inst_3_40(.clk(clk),.reset(reset),.i1(intermediate_reg_2[479]),.i2(intermediate_reg_2[478]),.o(intermediate_reg_3[239]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_41(.clk(clk),.reset(reset),.i1(intermediate_reg_2[477]),.i2(intermediate_reg_2[476]),.o(intermediate_reg_3[238]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_42(.clk(clk),.reset(reset),.i1(intermediate_reg_2[475]),.i2(intermediate_reg_2[474]),.o(intermediate_reg_3[237])); 
fsm fsm_inst_3_43(.clk(clk),.reset(reset),.i1(intermediate_reg_2[473]),.i2(intermediate_reg_2[472]),.o(intermediate_reg_3[236])); 
fsm fsm_inst_3_44(.clk(clk),.reset(reset),.i1(intermediate_reg_2[471]),.i2(intermediate_reg_2[470]),.o(intermediate_reg_3[235])); 
fsm fsm_inst_3_45(.clk(clk),.reset(reset),.i1(intermediate_reg_2[469]),.i2(intermediate_reg_2[468]),.o(intermediate_reg_3[234])); 
fsm fsm_inst_3_46(.clk(clk),.reset(reset),.i1(intermediate_reg_2[467]),.i2(intermediate_reg_2[466]),.o(intermediate_reg_3[233])); 
fsm fsm_inst_3_47(.clk(clk),.reset(reset),.i1(intermediate_reg_2[465]),.i2(intermediate_reg_2[464]),.o(intermediate_reg_3[232])); 
fsm fsm_inst_3_48(.clk(clk),.reset(reset),.i1(intermediate_reg_2[463]),.i2(intermediate_reg_2[462]),.o(intermediate_reg_3[231])); 
mux_module mux_module_inst_3_49(.clk(clk),.reset(reset),.i1(intermediate_reg_2[461]),.i2(intermediate_reg_2[460]),.o(intermediate_reg_3[230]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_50(.clk(clk),.reset(reset),.i1(intermediate_reg_2[459]),.i2(intermediate_reg_2[458]),.o(intermediate_reg_3[229]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_51(.clk(clk),.reset(reset),.i1(intermediate_reg_2[457]),.i2(intermediate_reg_2[456]),.o(intermediate_reg_3[228])); 
mux_module mux_module_inst_3_52(.clk(clk),.reset(reset),.i1(intermediate_reg_2[455]),.i2(intermediate_reg_2[454]),.o(intermediate_reg_3[227]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_53(.clk(clk),.reset(reset),.i1(intermediate_reg_2[453]),.i2(intermediate_reg_2[452]),.o(intermediate_reg_3[226])); 
mux_module mux_module_inst_3_54(.clk(clk),.reset(reset),.i1(intermediate_reg_2[451]),.i2(intermediate_reg_2[450]),.o(intermediate_reg_3[225]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_55(.clk(clk),.reset(reset),.i1(intermediate_reg_2[449]),.i2(intermediate_reg_2[448]),.o(intermediate_reg_3[224]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_56(.clk(clk),.reset(reset),.i1(intermediate_reg_2[447]),.i2(intermediate_reg_2[446]),.o(intermediate_reg_3[223])); 
fsm fsm_inst_3_57(.clk(clk),.reset(reset),.i1(intermediate_reg_2[445]),.i2(intermediate_reg_2[444]),.o(intermediate_reg_3[222])); 
mux_module mux_module_inst_3_58(.clk(clk),.reset(reset),.i1(intermediate_reg_2[443]),.i2(intermediate_reg_2[442]),.o(intermediate_reg_3[221]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_59(.clk(clk),.reset(reset),.i1(intermediate_reg_2[441]),.i2(intermediate_reg_2[440]),.o(intermediate_reg_3[220])); 
fsm fsm_inst_3_60(.clk(clk),.reset(reset),.i1(intermediate_reg_2[439]),.i2(intermediate_reg_2[438]),.o(intermediate_reg_3[219])); 
fsm fsm_inst_3_61(.clk(clk),.reset(reset),.i1(intermediate_reg_2[437]),.i2(intermediate_reg_2[436]),.o(intermediate_reg_3[218])); 
fsm fsm_inst_3_62(.clk(clk),.reset(reset),.i1(intermediate_reg_2[435]),.i2(intermediate_reg_2[434]),.o(intermediate_reg_3[217])); 
fsm fsm_inst_3_63(.clk(clk),.reset(reset),.i1(intermediate_reg_2[433]),.i2(intermediate_reg_2[432]),.o(intermediate_reg_3[216])); 
fsm fsm_inst_3_64(.clk(clk),.reset(reset),.i1(intermediate_reg_2[431]),.i2(intermediate_reg_2[430]),.o(intermediate_reg_3[215])); 
mux_module mux_module_inst_3_65(.clk(clk),.reset(reset),.i1(intermediate_reg_2[429]),.i2(intermediate_reg_2[428]),.o(intermediate_reg_3[214]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_66(.clk(clk),.reset(reset),.i1(intermediate_reg_2[427]),.i2(intermediate_reg_2[426]),.o(intermediate_reg_3[213]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_67(.clk(clk),.reset(reset),.i1(intermediate_reg_2[425]),.i2(intermediate_reg_2[424]),.o(intermediate_reg_3[212]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_68(.clk(clk),.reset(reset),.i1(intermediate_reg_2[423]),.i2(intermediate_reg_2[422]),.o(intermediate_reg_3[211]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_69(.clk(clk),.reset(reset),.i1(intermediate_reg_2[421]),.i2(intermediate_reg_2[420]),.o(intermediate_reg_3[210])); 
mux_module mux_module_inst_3_70(.clk(clk),.reset(reset),.i1(intermediate_reg_2[419]),.i2(intermediate_reg_2[418]),.o(intermediate_reg_3[209]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_71(.clk(clk),.reset(reset),.i1(intermediate_reg_2[417]),.i2(intermediate_reg_2[416]),.o(intermediate_reg_3[208])); 
fsm fsm_inst_3_72(.clk(clk),.reset(reset),.i1(intermediate_reg_2[415]),.i2(intermediate_reg_2[414]),.o(intermediate_reg_3[207])); 
mux_module mux_module_inst_3_73(.clk(clk),.reset(reset),.i1(intermediate_reg_2[413]),.i2(intermediate_reg_2[412]),.o(intermediate_reg_3[206]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_74(.clk(clk),.reset(reset),.i1(intermediate_reg_2[411]),.i2(intermediate_reg_2[410]),.o(intermediate_reg_3[205]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_75(.clk(clk),.reset(reset),.i1(intermediate_reg_2[409]),.i2(intermediate_reg_2[408]),.o(intermediate_reg_3[204])); 
mux_module mux_module_inst_3_76(.clk(clk),.reset(reset),.i1(intermediate_reg_2[407]),.i2(intermediate_reg_2[406]),.o(intermediate_reg_3[203]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_77(.clk(clk),.reset(reset),.i1(intermediate_reg_2[405]),.i2(intermediate_reg_2[404]),.o(intermediate_reg_3[202]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_78(.clk(clk),.reset(reset),.i1(intermediate_reg_2[403]),.i2(intermediate_reg_2[402]),.o(intermediate_reg_3[201]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_79(.clk(clk),.reset(reset),.i1(intermediate_reg_2[401]),.i2(intermediate_reg_2[400]),.o(intermediate_reg_3[200]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_80(.clk(clk),.reset(reset),.i1(intermediate_reg_2[399]),.i2(intermediate_reg_2[398]),.o(intermediate_reg_3[199]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_81(.clk(clk),.reset(reset),.i1(intermediate_reg_2[397]),.i2(intermediate_reg_2[396]),.o(intermediate_reg_3[198])); 
fsm fsm_inst_3_82(.clk(clk),.reset(reset),.i1(intermediate_reg_2[395]),.i2(intermediate_reg_2[394]),.o(intermediate_reg_3[197])); 
fsm fsm_inst_3_83(.clk(clk),.reset(reset),.i1(intermediate_reg_2[393]),.i2(intermediate_reg_2[392]),.o(intermediate_reg_3[196])); 
fsm fsm_inst_3_84(.clk(clk),.reset(reset),.i1(intermediate_reg_2[391]),.i2(intermediate_reg_2[390]),.o(intermediate_reg_3[195])); 
fsm fsm_inst_3_85(.clk(clk),.reset(reset),.i1(intermediate_reg_2[389]),.i2(intermediate_reg_2[388]),.o(intermediate_reg_3[194])); 
mux_module mux_module_inst_3_86(.clk(clk),.reset(reset),.i1(intermediate_reg_2[387]),.i2(intermediate_reg_2[386]),.o(intermediate_reg_3[193]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_87(.clk(clk),.reset(reset),.i1(intermediate_reg_2[385]),.i2(intermediate_reg_2[384]),.o(intermediate_reg_3[192])); 
fsm fsm_inst_3_88(.clk(clk),.reset(reset),.i1(intermediate_reg_2[383]),.i2(intermediate_reg_2[382]),.o(intermediate_reg_3[191])); 
fsm fsm_inst_3_89(.clk(clk),.reset(reset),.i1(intermediate_reg_2[381]),.i2(intermediate_reg_2[380]),.o(intermediate_reg_3[190])); 
fsm fsm_inst_3_90(.clk(clk),.reset(reset),.i1(intermediate_reg_2[379]),.i2(intermediate_reg_2[378]),.o(intermediate_reg_3[189])); 
mux_module mux_module_inst_3_91(.clk(clk),.reset(reset),.i1(intermediate_reg_2[377]),.i2(intermediate_reg_2[376]),.o(intermediate_reg_3[188]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_92(.clk(clk),.reset(reset),.i1(intermediate_reg_2[375]),.i2(intermediate_reg_2[374]),.o(intermediate_reg_3[187]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_93(.clk(clk),.reset(reset),.i1(intermediate_reg_2[373]),.i2(intermediate_reg_2[372]),.o(intermediate_reg_3[186]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_94(.clk(clk),.reset(reset),.i1(intermediate_reg_2[371]),.i2(intermediate_reg_2[370]),.o(intermediate_reg_3[185]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_95(.clk(clk),.reset(reset),.i1(intermediate_reg_2[369]),.i2(intermediate_reg_2[368]),.o(intermediate_reg_3[184]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_96(.clk(clk),.reset(reset),.i1(intermediate_reg_2[367]),.i2(intermediate_reg_2[366]),.o(intermediate_reg_3[183]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_97(.clk(clk),.reset(reset),.i1(intermediate_reg_2[365]),.i2(intermediate_reg_2[364]),.o(intermediate_reg_3[182]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_98(.clk(clk),.reset(reset),.i1(intermediate_reg_2[363]),.i2(intermediate_reg_2[362]),.o(intermediate_reg_3[181])); 
fsm fsm_inst_3_99(.clk(clk),.reset(reset),.i1(intermediate_reg_2[361]),.i2(intermediate_reg_2[360]),.o(intermediate_reg_3[180])); 
mux_module mux_module_inst_3_100(.clk(clk),.reset(reset),.i1(intermediate_reg_2[359]),.i2(intermediate_reg_2[358]),.o(intermediate_reg_3[179]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_101(.clk(clk),.reset(reset),.i1(intermediate_reg_2[357]),.i2(intermediate_reg_2[356]),.o(intermediate_reg_3[178]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_102(.clk(clk),.reset(reset),.i1(intermediate_reg_2[355]),.i2(intermediate_reg_2[354]),.o(intermediate_reg_3[177])); 
mux_module mux_module_inst_3_103(.clk(clk),.reset(reset),.i1(intermediate_reg_2[353]),.i2(intermediate_reg_2[352]),.o(intermediate_reg_3[176]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_104(.clk(clk),.reset(reset),.i1(intermediate_reg_2[351]),.i2(intermediate_reg_2[350]),.o(intermediate_reg_3[175]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_105(.clk(clk),.reset(reset),.i1(intermediate_reg_2[349]),.i2(intermediate_reg_2[348]),.o(intermediate_reg_3[174])); 
fsm fsm_inst_3_106(.clk(clk),.reset(reset),.i1(intermediate_reg_2[347]),.i2(intermediate_reg_2[346]),.o(intermediate_reg_3[173])); 
mux_module mux_module_inst_3_107(.clk(clk),.reset(reset),.i1(intermediate_reg_2[345]),.i2(intermediate_reg_2[344]),.o(intermediate_reg_3[172]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_108(.clk(clk),.reset(reset),.i1(intermediate_reg_2[343]),.i2(intermediate_reg_2[342]),.o(intermediate_reg_3[171]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_109(.clk(clk),.reset(reset),.i1(intermediate_reg_2[341]),.i2(intermediate_reg_2[340]),.o(intermediate_reg_3[170])); 
mux_module mux_module_inst_3_110(.clk(clk),.reset(reset),.i1(intermediate_reg_2[339]),.i2(intermediate_reg_2[338]),.o(intermediate_reg_3[169]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_111(.clk(clk),.reset(reset),.i1(intermediate_reg_2[337]),.i2(intermediate_reg_2[336]),.o(intermediate_reg_3[168])); 
mux_module mux_module_inst_3_112(.clk(clk),.reset(reset),.i1(intermediate_reg_2[335]),.i2(intermediate_reg_2[334]),.o(intermediate_reg_3[167]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_113(.clk(clk),.reset(reset),.i1(intermediate_reg_2[333]),.i2(intermediate_reg_2[332]),.o(intermediate_reg_3[166]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_114(.clk(clk),.reset(reset),.i1(intermediate_reg_2[331]),.i2(intermediate_reg_2[330]),.o(intermediate_reg_3[165])); 
fsm fsm_inst_3_115(.clk(clk),.reset(reset),.i1(intermediate_reg_2[329]),.i2(intermediate_reg_2[328]),.o(intermediate_reg_3[164])); 
fsm fsm_inst_3_116(.clk(clk),.reset(reset),.i1(intermediate_reg_2[327]),.i2(intermediate_reg_2[326]),.o(intermediate_reg_3[163])); 
fsm fsm_inst_3_117(.clk(clk),.reset(reset),.i1(intermediate_reg_2[325]),.i2(intermediate_reg_2[324]),.o(intermediate_reg_3[162])); 
fsm fsm_inst_3_118(.clk(clk),.reset(reset),.i1(intermediate_reg_2[323]),.i2(intermediate_reg_2[322]),.o(intermediate_reg_3[161])); 
mux_module mux_module_inst_3_119(.clk(clk),.reset(reset),.i1(intermediate_reg_2[321]),.i2(intermediate_reg_2[320]),.o(intermediate_reg_3[160]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_120(.clk(clk),.reset(reset),.i1(intermediate_reg_2[319]),.i2(intermediate_reg_2[318]),.o(intermediate_reg_3[159])); 
mux_module mux_module_inst_3_121(.clk(clk),.reset(reset),.i1(intermediate_reg_2[317]),.i2(intermediate_reg_2[316]),.o(intermediate_reg_3[158]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_122(.clk(clk),.reset(reset),.i1(intermediate_reg_2[315]),.i2(intermediate_reg_2[314]),.o(intermediate_reg_3[157]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_123(.clk(clk),.reset(reset),.i1(intermediate_reg_2[313]),.i2(intermediate_reg_2[312]),.o(intermediate_reg_3[156])); 
fsm fsm_inst_3_124(.clk(clk),.reset(reset),.i1(intermediate_reg_2[311]),.i2(intermediate_reg_2[310]),.o(intermediate_reg_3[155])); 
mux_module mux_module_inst_3_125(.clk(clk),.reset(reset),.i1(intermediate_reg_2[309]),.i2(intermediate_reg_2[308]),.o(intermediate_reg_3[154]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_126(.clk(clk),.reset(reset),.i1(intermediate_reg_2[307]),.i2(intermediate_reg_2[306]),.o(intermediate_reg_3[153])); 
mux_module mux_module_inst_3_127(.clk(clk),.reset(reset),.i1(intermediate_reg_2[305]),.i2(intermediate_reg_2[304]),.o(intermediate_reg_3[152]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_128(.clk(clk),.reset(reset),.i1(intermediate_reg_2[303]),.i2(intermediate_reg_2[302]),.o(intermediate_reg_3[151])); 
fsm fsm_inst_3_129(.clk(clk),.reset(reset),.i1(intermediate_reg_2[301]),.i2(intermediate_reg_2[300]),.o(intermediate_reg_3[150])); 
mux_module mux_module_inst_3_130(.clk(clk),.reset(reset),.i1(intermediate_reg_2[299]),.i2(intermediate_reg_2[298]),.o(intermediate_reg_3[149]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_131(.clk(clk),.reset(reset),.i1(intermediate_reg_2[297]),.i2(intermediate_reg_2[296]),.o(intermediate_reg_3[148])); 
mux_module mux_module_inst_3_132(.clk(clk),.reset(reset),.i1(intermediate_reg_2[295]),.i2(intermediate_reg_2[294]),.o(intermediate_reg_3[147]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_133(.clk(clk),.reset(reset),.i1(intermediate_reg_2[293]),.i2(intermediate_reg_2[292]),.o(intermediate_reg_3[146])); 
mux_module mux_module_inst_3_134(.clk(clk),.reset(reset),.i1(intermediate_reg_2[291]),.i2(intermediate_reg_2[290]),.o(intermediate_reg_3[145]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_135(.clk(clk),.reset(reset),.i1(intermediate_reg_2[289]),.i2(intermediate_reg_2[288]),.o(intermediate_reg_3[144]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_136(.clk(clk),.reset(reset),.i1(intermediate_reg_2[287]),.i2(intermediate_reg_2[286]),.o(intermediate_reg_3[143]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_137(.clk(clk),.reset(reset),.i1(intermediate_reg_2[285]),.i2(intermediate_reg_2[284]),.o(intermediate_reg_3[142]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_138(.clk(clk),.reset(reset),.i1(intermediate_reg_2[283]),.i2(intermediate_reg_2[282]),.o(intermediate_reg_3[141])); 
fsm fsm_inst_3_139(.clk(clk),.reset(reset),.i1(intermediate_reg_2[281]),.i2(intermediate_reg_2[280]),.o(intermediate_reg_3[140])); 
mux_module mux_module_inst_3_140(.clk(clk),.reset(reset),.i1(intermediate_reg_2[279]),.i2(intermediate_reg_2[278]),.o(intermediate_reg_3[139]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_141(.clk(clk),.reset(reset),.i1(intermediate_reg_2[277]),.i2(intermediate_reg_2[276]),.o(intermediate_reg_3[138]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_142(.clk(clk),.reset(reset),.i1(intermediate_reg_2[275]),.i2(intermediate_reg_2[274]),.o(intermediate_reg_3[137]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_143(.clk(clk),.reset(reset),.i1(intermediate_reg_2[273]),.i2(intermediate_reg_2[272]),.o(intermediate_reg_3[136]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_144(.clk(clk),.reset(reset),.i1(intermediate_reg_2[271]),.i2(intermediate_reg_2[270]),.o(intermediate_reg_3[135]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_145(.clk(clk),.reset(reset),.i1(intermediate_reg_2[269]),.i2(intermediate_reg_2[268]),.o(intermediate_reg_3[134]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_146(.clk(clk),.reset(reset),.i1(intermediate_reg_2[267]),.i2(intermediate_reg_2[266]),.o(intermediate_reg_3[133]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_147(.clk(clk),.reset(reset),.i1(intermediate_reg_2[265]),.i2(intermediate_reg_2[264]),.o(intermediate_reg_3[132]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_148(.clk(clk),.reset(reset),.i1(intermediate_reg_2[263]),.i2(intermediate_reg_2[262]),.o(intermediate_reg_3[131]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_149(.clk(clk),.reset(reset),.i1(intermediate_reg_2[261]),.i2(intermediate_reg_2[260]),.o(intermediate_reg_3[130])); 
mux_module mux_module_inst_3_150(.clk(clk),.reset(reset),.i1(intermediate_reg_2[259]),.i2(intermediate_reg_2[258]),.o(intermediate_reg_3[129]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_151(.clk(clk),.reset(reset),.i1(intermediate_reg_2[257]),.i2(intermediate_reg_2[256]),.o(intermediate_reg_3[128]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_152(.clk(clk),.reset(reset),.i1(intermediate_reg_2[255]),.i2(intermediate_reg_2[254]),.o(intermediate_reg_3[127]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_153(.clk(clk),.reset(reset),.i1(intermediate_reg_2[253]),.i2(intermediate_reg_2[252]),.o(intermediate_reg_3[126])); 
fsm fsm_inst_3_154(.clk(clk),.reset(reset),.i1(intermediate_reg_2[251]),.i2(intermediate_reg_2[250]),.o(intermediate_reg_3[125])); 
fsm fsm_inst_3_155(.clk(clk),.reset(reset),.i1(intermediate_reg_2[249]),.i2(intermediate_reg_2[248]),.o(intermediate_reg_3[124])); 
mux_module mux_module_inst_3_156(.clk(clk),.reset(reset),.i1(intermediate_reg_2[247]),.i2(intermediate_reg_2[246]),.o(intermediate_reg_3[123]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_157(.clk(clk),.reset(reset),.i1(intermediate_reg_2[245]),.i2(intermediate_reg_2[244]),.o(intermediate_reg_3[122])); 
mux_module mux_module_inst_3_158(.clk(clk),.reset(reset),.i1(intermediate_reg_2[243]),.i2(intermediate_reg_2[242]),.o(intermediate_reg_3[121]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_159(.clk(clk),.reset(reset),.i1(intermediate_reg_2[241]),.i2(intermediate_reg_2[240]),.o(intermediate_reg_3[120])); 
fsm fsm_inst_3_160(.clk(clk),.reset(reset),.i1(intermediate_reg_2[239]),.i2(intermediate_reg_2[238]),.o(intermediate_reg_3[119])); 
fsm fsm_inst_3_161(.clk(clk),.reset(reset),.i1(intermediate_reg_2[237]),.i2(intermediate_reg_2[236]),.o(intermediate_reg_3[118])); 
mux_module mux_module_inst_3_162(.clk(clk),.reset(reset),.i1(intermediate_reg_2[235]),.i2(intermediate_reg_2[234]),.o(intermediate_reg_3[117]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_163(.clk(clk),.reset(reset),.i1(intermediate_reg_2[233]),.i2(intermediate_reg_2[232]),.o(intermediate_reg_3[116]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_164(.clk(clk),.reset(reset),.i1(intermediate_reg_2[231]),.i2(intermediate_reg_2[230]),.o(intermediate_reg_3[115]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_165(.clk(clk),.reset(reset),.i1(intermediate_reg_2[229]),.i2(intermediate_reg_2[228]),.o(intermediate_reg_3[114])); 
mux_module mux_module_inst_3_166(.clk(clk),.reset(reset),.i1(intermediate_reg_2[227]),.i2(intermediate_reg_2[226]),.o(intermediate_reg_3[113]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_167(.clk(clk),.reset(reset),.i1(intermediate_reg_2[225]),.i2(intermediate_reg_2[224]),.o(intermediate_reg_3[112])); 
mux_module mux_module_inst_3_168(.clk(clk),.reset(reset),.i1(intermediate_reg_2[223]),.i2(intermediate_reg_2[222]),.o(intermediate_reg_3[111]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_169(.clk(clk),.reset(reset),.i1(intermediate_reg_2[221]),.i2(intermediate_reg_2[220]),.o(intermediate_reg_3[110]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_170(.clk(clk),.reset(reset),.i1(intermediate_reg_2[219]),.i2(intermediate_reg_2[218]),.o(intermediate_reg_3[109])); 
mux_module mux_module_inst_3_171(.clk(clk),.reset(reset),.i1(intermediate_reg_2[217]),.i2(intermediate_reg_2[216]),.o(intermediate_reg_3[108]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_172(.clk(clk),.reset(reset),.i1(intermediate_reg_2[215]),.i2(intermediate_reg_2[214]),.o(intermediate_reg_3[107])); 
mux_module mux_module_inst_3_173(.clk(clk),.reset(reset),.i1(intermediate_reg_2[213]),.i2(intermediate_reg_2[212]),.o(intermediate_reg_3[106]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_174(.clk(clk),.reset(reset),.i1(intermediate_reg_2[211]),.i2(intermediate_reg_2[210]),.o(intermediate_reg_3[105])); 
fsm fsm_inst_3_175(.clk(clk),.reset(reset),.i1(intermediate_reg_2[209]),.i2(intermediate_reg_2[208]),.o(intermediate_reg_3[104])); 
fsm fsm_inst_3_176(.clk(clk),.reset(reset),.i1(intermediate_reg_2[207]),.i2(intermediate_reg_2[206]),.o(intermediate_reg_3[103])); 
mux_module mux_module_inst_3_177(.clk(clk),.reset(reset),.i1(intermediate_reg_2[205]),.i2(intermediate_reg_2[204]),.o(intermediate_reg_3[102]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_178(.clk(clk),.reset(reset),.i1(intermediate_reg_2[203]),.i2(intermediate_reg_2[202]),.o(intermediate_reg_3[101]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_179(.clk(clk),.reset(reset),.i1(intermediate_reg_2[201]),.i2(intermediate_reg_2[200]),.o(intermediate_reg_3[100]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_180(.clk(clk),.reset(reset),.i1(intermediate_reg_2[199]),.i2(intermediate_reg_2[198]),.o(intermediate_reg_3[99]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_181(.clk(clk),.reset(reset),.i1(intermediate_reg_2[197]),.i2(intermediate_reg_2[196]),.o(intermediate_reg_3[98])); 
mux_module mux_module_inst_3_182(.clk(clk),.reset(reset),.i1(intermediate_reg_2[195]),.i2(intermediate_reg_2[194]),.o(intermediate_reg_3[97]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_183(.clk(clk),.reset(reset),.i1(intermediate_reg_2[193]),.i2(intermediate_reg_2[192]),.o(intermediate_reg_3[96])); 
fsm fsm_inst_3_184(.clk(clk),.reset(reset),.i1(intermediate_reg_2[191]),.i2(intermediate_reg_2[190]),.o(intermediate_reg_3[95])); 
fsm fsm_inst_3_185(.clk(clk),.reset(reset),.i1(intermediate_reg_2[189]),.i2(intermediate_reg_2[188]),.o(intermediate_reg_3[94])); 
fsm fsm_inst_3_186(.clk(clk),.reset(reset),.i1(intermediate_reg_2[187]),.i2(intermediate_reg_2[186]),.o(intermediate_reg_3[93])); 
fsm fsm_inst_3_187(.clk(clk),.reset(reset),.i1(intermediate_reg_2[185]),.i2(intermediate_reg_2[184]),.o(intermediate_reg_3[92])); 
fsm fsm_inst_3_188(.clk(clk),.reset(reset),.i1(intermediate_reg_2[183]),.i2(intermediate_reg_2[182]),.o(intermediate_reg_3[91])); 
mux_module mux_module_inst_3_189(.clk(clk),.reset(reset),.i1(intermediate_reg_2[181]),.i2(intermediate_reg_2[180]),.o(intermediate_reg_3[90]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_190(.clk(clk),.reset(reset),.i1(intermediate_reg_2[179]),.i2(intermediate_reg_2[178]),.o(intermediate_reg_3[89])); 
mux_module mux_module_inst_3_191(.clk(clk),.reset(reset),.i1(intermediate_reg_2[177]),.i2(intermediate_reg_2[176]),.o(intermediate_reg_3[88]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_192(.clk(clk),.reset(reset),.i1(intermediate_reg_2[175]),.i2(intermediate_reg_2[174]),.o(intermediate_reg_3[87]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_193(.clk(clk),.reset(reset),.i1(intermediate_reg_2[173]),.i2(intermediate_reg_2[172]),.o(intermediate_reg_3[86]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_194(.clk(clk),.reset(reset),.i1(intermediate_reg_2[171]),.i2(intermediate_reg_2[170]),.o(intermediate_reg_3[85]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_195(.clk(clk),.reset(reset),.i1(intermediate_reg_2[169]),.i2(intermediate_reg_2[168]),.o(intermediate_reg_3[84]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_196(.clk(clk),.reset(reset),.i1(intermediate_reg_2[167]),.i2(intermediate_reg_2[166]),.o(intermediate_reg_3[83])); 
mux_module mux_module_inst_3_197(.clk(clk),.reset(reset),.i1(intermediate_reg_2[165]),.i2(intermediate_reg_2[164]),.o(intermediate_reg_3[82]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_198(.clk(clk),.reset(reset),.i1(intermediate_reg_2[163]),.i2(intermediate_reg_2[162]),.o(intermediate_reg_3[81])); 
mux_module mux_module_inst_3_199(.clk(clk),.reset(reset),.i1(intermediate_reg_2[161]),.i2(intermediate_reg_2[160]),.o(intermediate_reg_3[80]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_200(.clk(clk),.reset(reset),.i1(intermediate_reg_2[159]),.i2(intermediate_reg_2[158]),.o(intermediate_reg_3[79]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_201(.clk(clk),.reset(reset),.i1(intermediate_reg_2[157]),.i2(intermediate_reg_2[156]),.o(intermediate_reg_3[78])); 
mux_module mux_module_inst_3_202(.clk(clk),.reset(reset),.i1(intermediate_reg_2[155]),.i2(intermediate_reg_2[154]),.o(intermediate_reg_3[77]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_203(.clk(clk),.reset(reset),.i1(intermediate_reg_2[153]),.i2(intermediate_reg_2[152]),.o(intermediate_reg_3[76]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_204(.clk(clk),.reset(reset),.i1(intermediate_reg_2[151]),.i2(intermediate_reg_2[150]),.o(intermediate_reg_3[75]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_205(.clk(clk),.reset(reset),.i1(intermediate_reg_2[149]),.i2(intermediate_reg_2[148]),.o(intermediate_reg_3[74]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_206(.clk(clk),.reset(reset),.i1(intermediate_reg_2[147]),.i2(intermediate_reg_2[146]),.o(intermediate_reg_3[73]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_207(.clk(clk),.reset(reset),.i1(intermediate_reg_2[145]),.i2(intermediate_reg_2[144]),.o(intermediate_reg_3[72]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_208(.clk(clk),.reset(reset),.i1(intermediate_reg_2[143]),.i2(intermediate_reg_2[142]),.o(intermediate_reg_3[71]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_209(.clk(clk),.reset(reset),.i1(intermediate_reg_2[141]),.i2(intermediate_reg_2[140]),.o(intermediate_reg_3[70]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_210(.clk(clk),.reset(reset),.i1(intermediate_reg_2[139]),.i2(intermediate_reg_2[138]),.o(intermediate_reg_3[69])); 
fsm fsm_inst_3_211(.clk(clk),.reset(reset),.i1(intermediate_reg_2[137]),.i2(intermediate_reg_2[136]),.o(intermediate_reg_3[68])); 
fsm fsm_inst_3_212(.clk(clk),.reset(reset),.i1(intermediate_reg_2[135]),.i2(intermediate_reg_2[134]),.o(intermediate_reg_3[67])); 
fsm fsm_inst_3_213(.clk(clk),.reset(reset),.i1(intermediate_reg_2[133]),.i2(intermediate_reg_2[132]),.o(intermediate_reg_3[66])); 
mux_module mux_module_inst_3_214(.clk(clk),.reset(reset),.i1(intermediate_reg_2[131]),.i2(intermediate_reg_2[130]),.o(intermediate_reg_3[65]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_215(.clk(clk),.reset(reset),.i1(intermediate_reg_2[129]),.i2(intermediate_reg_2[128]),.o(intermediate_reg_3[64])); 
fsm fsm_inst_3_216(.clk(clk),.reset(reset),.i1(intermediate_reg_2[127]),.i2(intermediate_reg_2[126]),.o(intermediate_reg_3[63])); 
mux_module mux_module_inst_3_217(.clk(clk),.reset(reset),.i1(intermediate_reg_2[125]),.i2(intermediate_reg_2[124]),.o(intermediate_reg_3[62]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_218(.clk(clk),.reset(reset),.i1(intermediate_reg_2[123]),.i2(intermediate_reg_2[122]),.o(intermediate_reg_3[61]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_219(.clk(clk),.reset(reset),.i1(intermediate_reg_2[121]),.i2(intermediate_reg_2[120]),.o(intermediate_reg_3[60])); 
mux_module mux_module_inst_3_220(.clk(clk),.reset(reset),.i1(intermediate_reg_2[119]),.i2(intermediate_reg_2[118]),.o(intermediate_reg_3[59]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_221(.clk(clk),.reset(reset),.i1(intermediate_reg_2[117]),.i2(intermediate_reg_2[116]),.o(intermediate_reg_3[58]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_222(.clk(clk),.reset(reset),.i1(intermediate_reg_2[115]),.i2(intermediate_reg_2[114]),.o(intermediate_reg_3[57])); 
fsm fsm_inst_3_223(.clk(clk),.reset(reset),.i1(intermediate_reg_2[113]),.i2(intermediate_reg_2[112]),.o(intermediate_reg_3[56])); 
mux_module mux_module_inst_3_224(.clk(clk),.reset(reset),.i1(intermediate_reg_2[111]),.i2(intermediate_reg_2[110]),.o(intermediate_reg_3[55]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_225(.clk(clk),.reset(reset),.i1(intermediate_reg_2[109]),.i2(intermediate_reg_2[108]),.o(intermediate_reg_3[54]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_226(.clk(clk),.reset(reset),.i1(intermediate_reg_2[107]),.i2(intermediate_reg_2[106]),.o(intermediate_reg_3[53])); 
mux_module mux_module_inst_3_227(.clk(clk),.reset(reset),.i1(intermediate_reg_2[105]),.i2(intermediate_reg_2[104]),.o(intermediate_reg_3[52]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_228(.clk(clk),.reset(reset),.i1(intermediate_reg_2[103]),.i2(intermediate_reg_2[102]),.o(intermediate_reg_3[51])); 
mux_module mux_module_inst_3_229(.clk(clk),.reset(reset),.i1(intermediate_reg_2[101]),.i2(intermediate_reg_2[100]),.o(intermediate_reg_3[50]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_230(.clk(clk),.reset(reset),.i1(intermediate_reg_2[99]),.i2(intermediate_reg_2[98]),.o(intermediate_reg_3[49]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_231(.clk(clk),.reset(reset),.i1(intermediate_reg_2[97]),.i2(intermediate_reg_2[96]),.o(intermediate_reg_3[48])); 
fsm fsm_inst_3_232(.clk(clk),.reset(reset),.i1(intermediate_reg_2[95]),.i2(intermediate_reg_2[94]),.o(intermediate_reg_3[47])); 
mux_module mux_module_inst_3_233(.clk(clk),.reset(reset),.i1(intermediate_reg_2[93]),.i2(intermediate_reg_2[92]),.o(intermediate_reg_3[46]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_234(.clk(clk),.reset(reset),.i1(intermediate_reg_2[91]),.i2(intermediate_reg_2[90]),.o(intermediate_reg_3[45])); 
mux_module mux_module_inst_3_235(.clk(clk),.reset(reset),.i1(intermediate_reg_2[89]),.i2(intermediate_reg_2[88]),.o(intermediate_reg_3[44]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_236(.clk(clk),.reset(reset),.i1(intermediate_reg_2[87]),.i2(intermediate_reg_2[86]),.o(intermediate_reg_3[43]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_237(.clk(clk),.reset(reset),.i1(intermediate_reg_2[85]),.i2(intermediate_reg_2[84]),.o(intermediate_reg_3[42])); 
fsm fsm_inst_3_238(.clk(clk),.reset(reset),.i1(intermediate_reg_2[83]),.i2(intermediate_reg_2[82]),.o(intermediate_reg_3[41])); 
fsm fsm_inst_3_239(.clk(clk),.reset(reset),.i1(intermediate_reg_2[81]),.i2(intermediate_reg_2[80]),.o(intermediate_reg_3[40])); 
fsm fsm_inst_3_240(.clk(clk),.reset(reset),.i1(intermediate_reg_2[79]),.i2(intermediate_reg_2[78]),.o(intermediate_reg_3[39])); 
fsm fsm_inst_3_241(.clk(clk),.reset(reset),.i1(intermediate_reg_2[77]),.i2(intermediate_reg_2[76]),.o(intermediate_reg_3[38])); 
fsm fsm_inst_3_242(.clk(clk),.reset(reset),.i1(intermediate_reg_2[75]),.i2(intermediate_reg_2[74]),.o(intermediate_reg_3[37])); 
fsm fsm_inst_3_243(.clk(clk),.reset(reset),.i1(intermediate_reg_2[73]),.i2(intermediate_reg_2[72]),.o(intermediate_reg_3[36])); 
mux_module mux_module_inst_3_244(.clk(clk),.reset(reset),.i1(intermediate_reg_2[71]),.i2(intermediate_reg_2[70]),.o(intermediate_reg_3[35]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_245(.clk(clk),.reset(reset),.i1(intermediate_reg_2[69]),.i2(intermediate_reg_2[68]),.o(intermediate_reg_3[34]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_246(.clk(clk),.reset(reset),.i1(intermediate_reg_2[67]),.i2(intermediate_reg_2[66]),.o(intermediate_reg_3[33]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_247(.clk(clk),.reset(reset),.i1(intermediate_reg_2[65]),.i2(intermediate_reg_2[64]),.o(intermediate_reg_3[32]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_248(.clk(clk),.reset(reset),.i1(intermediate_reg_2[63]),.i2(intermediate_reg_2[62]),.o(intermediate_reg_3[31])); 
fsm fsm_inst_3_249(.clk(clk),.reset(reset),.i1(intermediate_reg_2[61]),.i2(intermediate_reg_2[60]),.o(intermediate_reg_3[30])); 
fsm fsm_inst_3_250(.clk(clk),.reset(reset),.i1(intermediate_reg_2[59]),.i2(intermediate_reg_2[58]),.o(intermediate_reg_3[29])); 
fsm fsm_inst_3_251(.clk(clk),.reset(reset),.i1(intermediate_reg_2[57]),.i2(intermediate_reg_2[56]),.o(intermediate_reg_3[28])); 
mux_module mux_module_inst_3_252(.clk(clk),.reset(reset),.i1(intermediate_reg_2[55]),.i2(intermediate_reg_2[54]),.o(intermediate_reg_3[27]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_253(.clk(clk),.reset(reset),.i1(intermediate_reg_2[53]),.i2(intermediate_reg_2[52]),.o(intermediate_reg_3[26]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_254(.clk(clk),.reset(reset),.i1(intermediate_reg_2[51]),.i2(intermediate_reg_2[50]),.o(intermediate_reg_3[25])); 
mux_module mux_module_inst_3_255(.clk(clk),.reset(reset),.i1(intermediate_reg_2[49]),.i2(intermediate_reg_2[48]),.o(intermediate_reg_3[24]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_256(.clk(clk),.reset(reset),.i1(intermediate_reg_2[47]),.i2(intermediate_reg_2[46]),.o(intermediate_reg_3[23]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_257(.clk(clk),.reset(reset),.i1(intermediate_reg_2[45]),.i2(intermediate_reg_2[44]),.o(intermediate_reg_3[22])); 
fsm fsm_inst_3_258(.clk(clk),.reset(reset),.i1(intermediate_reg_2[43]),.i2(intermediate_reg_2[42]),.o(intermediate_reg_3[21])); 
fsm fsm_inst_3_259(.clk(clk),.reset(reset),.i1(intermediate_reg_2[41]),.i2(intermediate_reg_2[40]),.o(intermediate_reg_3[20])); 
mux_module mux_module_inst_3_260(.clk(clk),.reset(reset),.i1(intermediate_reg_2[39]),.i2(intermediate_reg_2[38]),.o(intermediate_reg_3[19]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_261(.clk(clk),.reset(reset),.i1(intermediate_reg_2[37]),.i2(intermediate_reg_2[36]),.o(intermediate_reg_3[18]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_262(.clk(clk),.reset(reset),.i1(intermediate_reg_2[35]),.i2(intermediate_reg_2[34]),.o(intermediate_reg_3[17]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_263(.clk(clk),.reset(reset),.i1(intermediate_reg_2[33]),.i2(intermediate_reg_2[32]),.o(intermediate_reg_3[16])); 
mux_module mux_module_inst_3_264(.clk(clk),.reset(reset),.i1(intermediate_reg_2[31]),.i2(intermediate_reg_2[30]),.o(intermediate_reg_3[15]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_265(.clk(clk),.reset(reset),.i1(intermediate_reg_2[29]),.i2(intermediate_reg_2[28]),.o(intermediate_reg_3[14]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_266(.clk(clk),.reset(reset),.i1(intermediate_reg_2[27]),.i2(intermediate_reg_2[26]),.o(intermediate_reg_3[13])); 
fsm fsm_inst_3_267(.clk(clk),.reset(reset),.i1(intermediate_reg_2[25]),.i2(intermediate_reg_2[24]),.o(intermediate_reg_3[12])); 
mux_module mux_module_inst_3_268(.clk(clk),.reset(reset),.i1(intermediate_reg_2[23]),.i2(intermediate_reg_2[22]),.o(intermediate_reg_3[11]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_269(.clk(clk),.reset(reset),.i1(intermediate_reg_2[21]),.i2(intermediate_reg_2[20]),.o(intermediate_reg_3[10]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_270(.clk(clk),.reset(reset),.i1(intermediate_reg_2[19]),.i2(intermediate_reg_2[18]),.o(intermediate_reg_3[9])); 
fsm fsm_inst_3_271(.clk(clk),.reset(reset),.i1(intermediate_reg_2[17]),.i2(intermediate_reg_2[16]),.o(intermediate_reg_3[8])); 
mux_module mux_module_inst_3_272(.clk(clk),.reset(reset),.i1(intermediate_reg_2[15]),.i2(intermediate_reg_2[14]),.o(intermediate_reg_3[7]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_273(.clk(clk),.reset(reset),.i1(intermediate_reg_2[13]),.i2(intermediate_reg_2[12]),.o(intermediate_reg_3[6]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_274(.clk(clk),.reset(reset),.i1(intermediate_reg_2[11]),.i2(intermediate_reg_2[10]),.o(intermediate_reg_3[5]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_275(.clk(clk),.reset(reset),.i1(intermediate_reg_2[9]),.i2(intermediate_reg_2[8]),.o(intermediate_reg_3[4]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_276(.clk(clk),.reset(reset),.i1(intermediate_reg_2[7]),.i2(intermediate_reg_2[6]),.o(intermediate_reg_3[3]),.sel(intermediate_reg_2[0])); 
mux_module mux_module_inst_3_277(.clk(clk),.reset(reset),.i1(intermediate_reg_2[5]),.i2(intermediate_reg_2[4]),.o(intermediate_reg_3[2]),.sel(intermediate_reg_2[0])); 
fsm fsm_inst_3_278(.clk(clk),.reset(reset),.i1(intermediate_reg_2[3]),.i2(intermediate_reg_2[2]),.o(intermediate_reg_3[1])); 
fsm fsm_inst_3_279(.clk(clk),.reset(reset),.i1(intermediate_reg_2[1]),.i2(intermediate_reg_2[0]),.o(intermediate_reg_3[0])); 
always@(posedge clk) begin 
outp [279:0] <= intermediate_reg_3; 
outp[527:280] <= intermediate_reg_3[247:0] ; 
end 
endmodule 
 

module interface_26(input reg [5359:0] inp, output reg [4319:0] outp, input clk, input reset);
reg [5359:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [2679:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5359]),.i2(intermediate_reg_0[5358]),.o(intermediate_reg_1[2679]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5357]),.i2(intermediate_reg_0[5356]),.o(intermediate_reg_1[2678]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5355]),.i2(intermediate_reg_0[5354]),.o(intermediate_reg_1[2677]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5353]),.i2(intermediate_reg_0[5352]),.o(intermediate_reg_1[2676])); 
fsm fsm_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5351]),.i2(intermediate_reg_0[5350]),.o(intermediate_reg_1[2675])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5349]),.i2(intermediate_reg_0[5348]),.o(intermediate_reg_1[2674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5347]),.i2(intermediate_reg_0[5346]),.o(intermediate_reg_1[2673]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5345]),.i2(intermediate_reg_0[5344]),.o(intermediate_reg_1[2672]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5343]),.i2(intermediate_reg_0[5342]),.o(intermediate_reg_1[2671])); 
fsm fsm_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5341]),.i2(intermediate_reg_0[5340]),.o(intermediate_reg_1[2670])); 
fsm fsm_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5339]),.i2(intermediate_reg_0[5338]),.o(intermediate_reg_1[2669])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5337]),.i2(intermediate_reg_0[5336]),.o(intermediate_reg_1[2668])); 
fsm fsm_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5335]),.i2(intermediate_reg_0[5334]),.o(intermediate_reg_1[2667])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5333]),.i2(intermediate_reg_0[5332]),.o(intermediate_reg_1[2666]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5331]),.i2(intermediate_reg_0[5330]),.o(intermediate_reg_1[2665])); 
fsm fsm_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5329]),.i2(intermediate_reg_0[5328]),.o(intermediate_reg_1[2664])); 
mux_module mux_module_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5327]),.i2(intermediate_reg_0[5326]),.o(intermediate_reg_1[2663]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5325]),.i2(intermediate_reg_0[5324]),.o(intermediate_reg_1[2662]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5323]),.i2(intermediate_reg_0[5322]),.o(intermediate_reg_1[2661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5321]),.i2(intermediate_reg_0[5320]),.o(intermediate_reg_1[2660]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5319]),.i2(intermediate_reg_0[5318]),.o(intermediate_reg_1[2659]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5317]),.i2(intermediate_reg_0[5316]),.o(intermediate_reg_1[2658])); 
fsm fsm_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5315]),.i2(intermediate_reg_0[5314]),.o(intermediate_reg_1[2657])); 
mux_module mux_module_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5313]),.i2(intermediate_reg_0[5312]),.o(intermediate_reg_1[2656]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5311]),.i2(intermediate_reg_0[5310]),.o(intermediate_reg_1[2655]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5309]),.i2(intermediate_reg_0[5308]),.o(intermediate_reg_1[2654])); 
mux_module mux_module_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5307]),.i2(intermediate_reg_0[5306]),.o(intermediate_reg_1[2653]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5305]),.i2(intermediate_reg_0[5304]),.o(intermediate_reg_1[2652]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5303]),.i2(intermediate_reg_0[5302]),.o(intermediate_reg_1[2651])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5301]),.i2(intermediate_reg_0[5300]),.o(intermediate_reg_1[2650]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5299]),.i2(intermediate_reg_0[5298]),.o(intermediate_reg_1[2649])); 
mux_module mux_module_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5297]),.i2(intermediate_reg_0[5296]),.o(intermediate_reg_1[2648]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5295]),.i2(intermediate_reg_0[5294]),.o(intermediate_reg_1[2647])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5293]),.i2(intermediate_reg_0[5292]),.o(intermediate_reg_1[2646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5291]),.i2(intermediate_reg_0[5290]),.o(intermediate_reg_1[2645]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5289]),.i2(intermediate_reg_0[5288]),.o(intermediate_reg_1[2644])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5287]),.i2(intermediate_reg_0[5286]),.o(intermediate_reg_1[2643]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5285]),.i2(intermediate_reg_0[5284]),.o(intermediate_reg_1[2642])); 
fsm fsm_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5283]),.i2(intermediate_reg_0[5282]),.o(intermediate_reg_1[2641])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5281]),.i2(intermediate_reg_0[5280]),.o(intermediate_reg_1[2640]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5279]),.i2(intermediate_reg_0[5278]),.o(intermediate_reg_1[2639])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5277]),.i2(intermediate_reg_0[5276]),.o(intermediate_reg_1[2638])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5275]),.i2(intermediate_reg_0[5274]),.o(intermediate_reg_1[2637]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5273]),.i2(intermediate_reg_0[5272]),.o(intermediate_reg_1[2636])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5271]),.i2(intermediate_reg_0[5270]),.o(intermediate_reg_1[2635]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5269]),.i2(intermediate_reg_0[5268]),.o(intermediate_reg_1[2634]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5267]),.i2(intermediate_reg_0[5266]),.o(intermediate_reg_1[2633]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5265]),.i2(intermediate_reg_0[5264]),.o(intermediate_reg_1[2632])); 
fsm fsm_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5263]),.i2(intermediate_reg_0[5262]),.o(intermediate_reg_1[2631])); 
fsm fsm_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5261]),.i2(intermediate_reg_0[5260]),.o(intermediate_reg_1[2630])); 
fsm fsm_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5259]),.i2(intermediate_reg_0[5258]),.o(intermediate_reg_1[2629])); 
fsm fsm_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5257]),.i2(intermediate_reg_0[5256]),.o(intermediate_reg_1[2628])); 
mux_module mux_module_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5255]),.i2(intermediate_reg_0[5254]),.o(intermediate_reg_1[2627]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5253]),.i2(intermediate_reg_0[5252]),.o(intermediate_reg_1[2626])); 
fsm fsm_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5251]),.i2(intermediate_reg_0[5250]),.o(intermediate_reg_1[2625])); 
fsm fsm_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5249]),.i2(intermediate_reg_0[5248]),.o(intermediate_reg_1[2624])); 
mux_module mux_module_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5247]),.i2(intermediate_reg_0[5246]),.o(intermediate_reg_1[2623]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5245]),.i2(intermediate_reg_0[5244]),.o(intermediate_reg_1[2622]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5243]),.i2(intermediate_reg_0[5242]),.o(intermediate_reg_1[2621])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5241]),.i2(intermediate_reg_0[5240]),.o(intermediate_reg_1[2620]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5239]),.i2(intermediate_reg_0[5238]),.o(intermediate_reg_1[2619])); 
mux_module mux_module_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5237]),.i2(intermediate_reg_0[5236]),.o(intermediate_reg_1[2618]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5235]),.i2(intermediate_reg_0[5234]),.o(intermediate_reg_1[2617])); 
fsm fsm_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5233]),.i2(intermediate_reg_0[5232]),.o(intermediate_reg_1[2616])); 
fsm fsm_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5231]),.i2(intermediate_reg_0[5230]),.o(intermediate_reg_1[2615])); 
mux_module mux_module_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5229]),.i2(intermediate_reg_0[5228]),.o(intermediate_reg_1[2614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5227]),.i2(intermediate_reg_0[5226]),.o(intermediate_reg_1[2613]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5225]),.i2(intermediate_reg_0[5224]),.o(intermediate_reg_1[2612]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5223]),.i2(intermediate_reg_0[5222]),.o(intermediate_reg_1[2611])); 
mux_module mux_module_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5221]),.i2(intermediate_reg_0[5220]),.o(intermediate_reg_1[2610]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5219]),.i2(intermediate_reg_0[5218]),.o(intermediate_reg_1[2609])); 
fsm fsm_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5217]),.i2(intermediate_reg_0[5216]),.o(intermediate_reg_1[2608])); 
fsm fsm_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5215]),.i2(intermediate_reg_0[5214]),.o(intermediate_reg_1[2607])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5213]),.i2(intermediate_reg_0[5212]),.o(intermediate_reg_1[2606]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5211]),.i2(intermediate_reg_0[5210]),.o(intermediate_reg_1[2605])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5209]),.i2(intermediate_reg_0[5208]),.o(intermediate_reg_1[2604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5207]),.i2(intermediate_reg_0[5206]),.o(intermediate_reg_1[2603]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5205]),.i2(intermediate_reg_0[5204]),.o(intermediate_reg_1[2602]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5203]),.i2(intermediate_reg_0[5202]),.o(intermediate_reg_1[2601])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5201]),.i2(intermediate_reg_0[5200]),.o(intermediate_reg_1[2600])); 
mux_module mux_module_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5199]),.i2(intermediate_reg_0[5198]),.o(intermediate_reg_1[2599]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5197]),.i2(intermediate_reg_0[5196]),.o(intermediate_reg_1[2598])); 
fsm fsm_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5195]),.i2(intermediate_reg_0[5194]),.o(intermediate_reg_1[2597])); 
fsm fsm_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5193]),.i2(intermediate_reg_0[5192]),.o(intermediate_reg_1[2596])); 
fsm fsm_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5191]),.i2(intermediate_reg_0[5190]),.o(intermediate_reg_1[2595])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5189]),.i2(intermediate_reg_0[5188]),.o(intermediate_reg_1[2594]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5187]),.i2(intermediate_reg_0[5186]),.o(intermediate_reg_1[2593]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5185]),.i2(intermediate_reg_0[5184]),.o(intermediate_reg_1[2592])); 
fsm fsm_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5183]),.i2(intermediate_reg_0[5182]),.o(intermediate_reg_1[2591])); 
fsm fsm_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5181]),.i2(intermediate_reg_0[5180]),.o(intermediate_reg_1[2590])); 
mux_module mux_module_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5179]),.i2(intermediate_reg_0[5178]),.o(intermediate_reg_1[2589]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5177]),.i2(intermediate_reg_0[5176]),.o(intermediate_reg_1[2588])); 
fsm fsm_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5175]),.i2(intermediate_reg_0[5174]),.o(intermediate_reg_1[2587])); 
fsm fsm_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5173]),.i2(intermediate_reg_0[5172]),.o(intermediate_reg_1[2586])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5171]),.i2(intermediate_reg_0[5170]),.o(intermediate_reg_1[2585]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5169]),.i2(intermediate_reg_0[5168]),.o(intermediate_reg_1[2584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5167]),.i2(intermediate_reg_0[5166]),.o(intermediate_reg_1[2583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5165]),.i2(intermediate_reg_0[5164]),.o(intermediate_reg_1[2582]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5163]),.i2(intermediate_reg_0[5162]),.o(intermediate_reg_1[2581]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5161]),.i2(intermediate_reg_0[5160]),.o(intermediate_reg_1[2580]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5159]),.i2(intermediate_reg_0[5158]),.o(intermediate_reg_1[2579])); 
fsm fsm_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5157]),.i2(intermediate_reg_0[5156]),.o(intermediate_reg_1[2578])); 
fsm fsm_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5155]),.i2(intermediate_reg_0[5154]),.o(intermediate_reg_1[2577])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5153]),.i2(intermediate_reg_0[5152]),.o(intermediate_reg_1[2576]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5151]),.i2(intermediate_reg_0[5150]),.o(intermediate_reg_1[2575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5149]),.i2(intermediate_reg_0[5148]),.o(intermediate_reg_1[2574]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5147]),.i2(intermediate_reg_0[5146]),.o(intermediate_reg_1[2573])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5145]),.i2(intermediate_reg_0[5144]),.o(intermediate_reg_1[2572]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5143]),.i2(intermediate_reg_0[5142]),.o(intermediate_reg_1[2571])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5141]),.i2(intermediate_reg_0[5140]),.o(intermediate_reg_1[2570]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5139]),.i2(intermediate_reg_0[5138]),.o(intermediate_reg_1[2569]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5137]),.i2(intermediate_reg_0[5136]),.o(intermediate_reg_1[2568]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5135]),.i2(intermediate_reg_0[5134]),.o(intermediate_reg_1[2567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5133]),.i2(intermediate_reg_0[5132]),.o(intermediate_reg_1[2566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5131]),.i2(intermediate_reg_0[5130]),.o(intermediate_reg_1[2565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5129]),.i2(intermediate_reg_0[5128]),.o(intermediate_reg_1[2564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5127]),.i2(intermediate_reg_0[5126]),.o(intermediate_reg_1[2563]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5125]),.i2(intermediate_reg_0[5124]),.o(intermediate_reg_1[2562])); 
mux_module mux_module_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5123]),.i2(intermediate_reg_0[5122]),.o(intermediate_reg_1[2561]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5121]),.i2(intermediate_reg_0[5120]),.o(intermediate_reg_1[2560]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5119]),.i2(intermediate_reg_0[5118]),.o(intermediate_reg_1[2559]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5117]),.i2(intermediate_reg_0[5116]),.o(intermediate_reg_1[2558])); 
mux_module mux_module_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5115]),.i2(intermediate_reg_0[5114]),.o(intermediate_reg_1[2557]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5113]),.i2(intermediate_reg_0[5112]),.o(intermediate_reg_1[2556])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5111]),.i2(intermediate_reg_0[5110]),.o(intermediate_reg_1[2555]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5109]),.i2(intermediate_reg_0[5108]),.o(intermediate_reg_1[2554])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5107]),.i2(intermediate_reg_0[5106]),.o(intermediate_reg_1[2553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5105]),.i2(intermediate_reg_0[5104]),.o(intermediate_reg_1[2552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5103]),.i2(intermediate_reg_0[5102]),.o(intermediate_reg_1[2551]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5101]),.i2(intermediate_reg_0[5100]),.o(intermediate_reg_1[2550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5099]),.i2(intermediate_reg_0[5098]),.o(intermediate_reg_1[2549]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5097]),.i2(intermediate_reg_0[5096]),.o(intermediate_reg_1[2548])); 
fsm fsm_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5095]),.i2(intermediate_reg_0[5094]),.o(intermediate_reg_1[2547])); 
mux_module mux_module_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5093]),.i2(intermediate_reg_0[5092]),.o(intermediate_reg_1[2546]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5091]),.i2(intermediate_reg_0[5090]),.o(intermediate_reg_1[2545])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5089]),.i2(intermediate_reg_0[5088]),.o(intermediate_reg_1[2544]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5087]),.i2(intermediate_reg_0[5086]),.o(intermediate_reg_1[2543])); 
fsm fsm_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5085]),.i2(intermediate_reg_0[5084]),.o(intermediate_reg_1[2542])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5083]),.i2(intermediate_reg_0[5082]),.o(intermediate_reg_1[2541]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5081]),.i2(intermediate_reg_0[5080]),.o(intermediate_reg_1[2540])); 
mux_module mux_module_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5079]),.i2(intermediate_reg_0[5078]),.o(intermediate_reg_1[2539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5077]),.i2(intermediate_reg_0[5076]),.o(intermediate_reg_1[2538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5075]),.i2(intermediate_reg_0[5074]),.o(intermediate_reg_1[2537]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5073]),.i2(intermediate_reg_0[5072]),.o(intermediate_reg_1[2536])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5071]),.i2(intermediate_reg_0[5070]),.o(intermediate_reg_1[2535]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5069]),.i2(intermediate_reg_0[5068]),.o(intermediate_reg_1[2534]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5067]),.i2(intermediate_reg_0[5066]),.o(intermediate_reg_1[2533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5065]),.i2(intermediate_reg_0[5064]),.o(intermediate_reg_1[2532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5063]),.i2(intermediate_reg_0[5062]),.o(intermediate_reg_1[2531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5061]),.i2(intermediate_reg_0[5060]),.o(intermediate_reg_1[2530]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5059]),.i2(intermediate_reg_0[5058]),.o(intermediate_reg_1[2529]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5057]),.i2(intermediate_reg_0[5056]),.o(intermediate_reg_1[2528])); 
mux_module mux_module_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5055]),.i2(intermediate_reg_0[5054]),.o(intermediate_reg_1[2527]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5053]),.i2(intermediate_reg_0[5052]),.o(intermediate_reg_1[2526])); 
fsm fsm_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5051]),.i2(intermediate_reg_0[5050]),.o(intermediate_reg_1[2525])); 
mux_module mux_module_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5049]),.i2(intermediate_reg_0[5048]),.o(intermediate_reg_1[2524]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5047]),.i2(intermediate_reg_0[5046]),.o(intermediate_reg_1[2523])); 
fsm fsm_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5045]),.i2(intermediate_reg_0[5044]),.o(intermediate_reg_1[2522])); 
fsm fsm_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5043]),.i2(intermediate_reg_0[5042]),.o(intermediate_reg_1[2521])); 
fsm fsm_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5041]),.i2(intermediate_reg_0[5040]),.o(intermediate_reg_1[2520])); 
fsm fsm_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5039]),.i2(intermediate_reg_0[5038]),.o(intermediate_reg_1[2519])); 
mux_module mux_module_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5037]),.i2(intermediate_reg_0[5036]),.o(intermediate_reg_1[2518]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5035]),.i2(intermediate_reg_0[5034]),.o(intermediate_reg_1[2517])); 
mux_module mux_module_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5033]),.i2(intermediate_reg_0[5032]),.o(intermediate_reg_1[2516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5031]),.i2(intermediate_reg_0[5030]),.o(intermediate_reg_1[2515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5029]),.i2(intermediate_reg_0[5028]),.o(intermediate_reg_1[2514]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5027]),.i2(intermediate_reg_0[5026]),.o(intermediate_reg_1[2513])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5025]),.i2(intermediate_reg_0[5024]),.o(intermediate_reg_1[2512]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5023]),.i2(intermediate_reg_0[5022]),.o(intermediate_reg_1[2511])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5021]),.i2(intermediate_reg_0[5020]),.o(intermediate_reg_1[2510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5019]),.i2(intermediate_reg_0[5018]),.o(intermediate_reg_1[2509]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5017]),.i2(intermediate_reg_0[5016]),.o(intermediate_reg_1[2508])); 
mux_module mux_module_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5015]),.i2(intermediate_reg_0[5014]),.o(intermediate_reg_1[2507]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5013]),.i2(intermediate_reg_0[5012]),.o(intermediate_reg_1[2506]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5011]),.i2(intermediate_reg_0[5010]),.o(intermediate_reg_1[2505]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5009]),.i2(intermediate_reg_0[5008]),.o(intermediate_reg_1[2504]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5007]),.i2(intermediate_reg_0[5006]),.o(intermediate_reg_1[2503])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5005]),.i2(intermediate_reg_0[5004]),.o(intermediate_reg_1[2502]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5003]),.i2(intermediate_reg_0[5002]),.o(intermediate_reg_1[2501])); 
mux_module mux_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5001]),.i2(intermediate_reg_0[5000]),.o(intermediate_reg_1[2500]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4999]),.i2(intermediate_reg_0[4998]),.o(intermediate_reg_1[2499])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4997]),.i2(intermediate_reg_0[4996]),.o(intermediate_reg_1[2498]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4995]),.i2(intermediate_reg_0[4994]),.o(intermediate_reg_1[2497]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4993]),.i2(intermediate_reg_0[4992]),.o(intermediate_reg_1[2496])); 
mux_module mux_module_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4991]),.i2(intermediate_reg_0[4990]),.o(intermediate_reg_1[2495]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4989]),.i2(intermediate_reg_0[4988]),.o(intermediate_reg_1[2494]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4987]),.i2(intermediate_reg_0[4986]),.o(intermediate_reg_1[2493])); 
fsm fsm_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4985]),.i2(intermediate_reg_0[4984]),.o(intermediate_reg_1[2492])); 
fsm fsm_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4983]),.i2(intermediate_reg_0[4982]),.o(intermediate_reg_1[2491])); 
mux_module mux_module_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4981]),.i2(intermediate_reg_0[4980]),.o(intermediate_reg_1[2490]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4979]),.i2(intermediate_reg_0[4978]),.o(intermediate_reg_1[2489]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4977]),.i2(intermediate_reg_0[4976]),.o(intermediate_reg_1[2488])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4975]),.i2(intermediate_reg_0[4974]),.o(intermediate_reg_1[2487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4973]),.i2(intermediate_reg_0[4972]),.o(intermediate_reg_1[2486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4971]),.i2(intermediate_reg_0[4970]),.o(intermediate_reg_1[2485]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4969]),.i2(intermediate_reg_0[4968]),.o(intermediate_reg_1[2484])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4967]),.i2(intermediate_reg_0[4966]),.o(intermediate_reg_1[2483])); 
fsm fsm_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4965]),.i2(intermediate_reg_0[4964]),.o(intermediate_reg_1[2482])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4963]),.i2(intermediate_reg_0[4962]),.o(intermediate_reg_1[2481]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4961]),.i2(intermediate_reg_0[4960]),.o(intermediate_reg_1[2480]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4959]),.i2(intermediate_reg_0[4958]),.o(intermediate_reg_1[2479])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4957]),.i2(intermediate_reg_0[4956]),.o(intermediate_reg_1[2478])); 
fsm fsm_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4955]),.i2(intermediate_reg_0[4954]),.o(intermediate_reg_1[2477])); 
fsm fsm_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4953]),.i2(intermediate_reg_0[4952]),.o(intermediate_reg_1[2476])); 
fsm fsm_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4951]),.i2(intermediate_reg_0[4950]),.o(intermediate_reg_1[2475])); 
mux_module mux_module_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4949]),.i2(intermediate_reg_0[4948]),.o(intermediate_reg_1[2474]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4947]),.i2(intermediate_reg_0[4946]),.o(intermediate_reg_1[2473]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4945]),.i2(intermediate_reg_0[4944]),.o(intermediate_reg_1[2472])); 
mux_module mux_module_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4943]),.i2(intermediate_reg_0[4942]),.o(intermediate_reg_1[2471]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4941]),.i2(intermediate_reg_0[4940]),.o(intermediate_reg_1[2470])); 
fsm fsm_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4939]),.i2(intermediate_reg_0[4938]),.o(intermediate_reg_1[2469])); 
fsm fsm_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4937]),.i2(intermediate_reg_0[4936]),.o(intermediate_reg_1[2468])); 
fsm fsm_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4935]),.i2(intermediate_reg_0[4934]),.o(intermediate_reg_1[2467])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4933]),.i2(intermediate_reg_0[4932]),.o(intermediate_reg_1[2466]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4931]),.i2(intermediate_reg_0[4930]),.o(intermediate_reg_1[2465])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4929]),.i2(intermediate_reg_0[4928]),.o(intermediate_reg_1[2464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4927]),.i2(intermediate_reg_0[4926]),.o(intermediate_reg_1[2463]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4925]),.i2(intermediate_reg_0[4924]),.o(intermediate_reg_1[2462])); 
mux_module mux_module_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4923]),.i2(intermediate_reg_0[4922]),.o(intermediate_reg_1[2461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4921]),.i2(intermediate_reg_0[4920]),.o(intermediate_reg_1[2460]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4919]),.i2(intermediate_reg_0[4918]),.o(intermediate_reg_1[2459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4917]),.i2(intermediate_reg_0[4916]),.o(intermediate_reg_1[2458]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4915]),.i2(intermediate_reg_0[4914]),.o(intermediate_reg_1[2457]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4913]),.i2(intermediate_reg_0[4912]),.o(intermediate_reg_1[2456])); 
mux_module mux_module_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4911]),.i2(intermediate_reg_0[4910]),.o(intermediate_reg_1[2455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4909]),.i2(intermediate_reg_0[4908]),.o(intermediate_reg_1[2454]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4907]),.i2(intermediate_reg_0[4906]),.o(intermediate_reg_1[2453])); 
fsm fsm_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4905]),.i2(intermediate_reg_0[4904]),.o(intermediate_reg_1[2452])); 
fsm fsm_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4903]),.i2(intermediate_reg_0[4902]),.o(intermediate_reg_1[2451])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4901]),.i2(intermediate_reg_0[4900]),.o(intermediate_reg_1[2450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4899]),.i2(intermediate_reg_0[4898]),.o(intermediate_reg_1[2449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4897]),.i2(intermediate_reg_0[4896]),.o(intermediate_reg_1[2448])); 
fsm fsm_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4895]),.i2(intermediate_reg_0[4894]),.o(intermediate_reg_1[2447])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4893]),.i2(intermediate_reg_0[4892]),.o(intermediate_reg_1[2446]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4891]),.i2(intermediate_reg_0[4890]),.o(intermediate_reg_1[2445])); 
fsm fsm_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4889]),.i2(intermediate_reg_0[4888]),.o(intermediate_reg_1[2444])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4887]),.i2(intermediate_reg_0[4886]),.o(intermediate_reg_1[2443])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4885]),.i2(intermediate_reg_0[4884]),.o(intermediate_reg_1[2442])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4883]),.i2(intermediate_reg_0[4882]),.o(intermediate_reg_1[2441]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4881]),.i2(intermediate_reg_0[4880]),.o(intermediate_reg_1[2440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4879]),.i2(intermediate_reg_0[4878]),.o(intermediate_reg_1[2439]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4877]),.i2(intermediate_reg_0[4876]),.o(intermediate_reg_1[2438]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4875]),.i2(intermediate_reg_0[4874]),.o(intermediate_reg_1[2437])); 
fsm fsm_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4873]),.i2(intermediate_reg_0[4872]),.o(intermediate_reg_1[2436])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4871]),.i2(intermediate_reg_0[4870]),.o(intermediate_reg_1[2435]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4869]),.i2(intermediate_reg_0[4868]),.o(intermediate_reg_1[2434]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4867]),.i2(intermediate_reg_0[4866]),.o(intermediate_reg_1[2433])); 
fsm fsm_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4865]),.i2(intermediate_reg_0[4864]),.o(intermediate_reg_1[2432])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4863]),.i2(intermediate_reg_0[4862]),.o(intermediate_reg_1[2431]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4861]),.i2(intermediate_reg_0[4860]),.o(intermediate_reg_1[2430])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4859]),.i2(intermediate_reg_0[4858]),.o(intermediate_reg_1[2429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4857]),.i2(intermediate_reg_0[4856]),.o(intermediate_reg_1[2428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4855]),.i2(intermediate_reg_0[4854]),.o(intermediate_reg_1[2427]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4853]),.i2(intermediate_reg_0[4852]),.o(intermediate_reg_1[2426])); 
fsm fsm_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4851]),.i2(intermediate_reg_0[4850]),.o(intermediate_reg_1[2425])); 
fsm fsm_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4849]),.i2(intermediate_reg_0[4848]),.o(intermediate_reg_1[2424])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4847]),.i2(intermediate_reg_0[4846]),.o(intermediate_reg_1[2423])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4845]),.i2(intermediate_reg_0[4844]),.o(intermediate_reg_1[2422]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4843]),.i2(intermediate_reg_0[4842]),.o(intermediate_reg_1[2421])); 
fsm fsm_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4841]),.i2(intermediate_reg_0[4840]),.o(intermediate_reg_1[2420])); 
fsm fsm_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4839]),.i2(intermediate_reg_0[4838]),.o(intermediate_reg_1[2419])); 
mux_module mux_module_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4837]),.i2(intermediate_reg_0[4836]),.o(intermediate_reg_1[2418]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4835]),.i2(intermediate_reg_0[4834]),.o(intermediate_reg_1[2417]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4833]),.i2(intermediate_reg_0[4832]),.o(intermediate_reg_1[2416])); 
mux_module mux_module_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4831]),.i2(intermediate_reg_0[4830]),.o(intermediate_reg_1[2415]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4829]),.i2(intermediate_reg_0[4828]),.o(intermediate_reg_1[2414]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4827]),.i2(intermediate_reg_0[4826]),.o(intermediate_reg_1[2413])); 
fsm fsm_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4825]),.i2(intermediate_reg_0[4824]),.o(intermediate_reg_1[2412])); 
mux_module mux_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4823]),.i2(intermediate_reg_0[4822]),.o(intermediate_reg_1[2411]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4821]),.i2(intermediate_reg_0[4820]),.o(intermediate_reg_1[2410]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4819]),.i2(intermediate_reg_0[4818]),.o(intermediate_reg_1[2409]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4817]),.i2(intermediate_reg_0[4816]),.o(intermediate_reg_1[2408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4815]),.i2(intermediate_reg_0[4814]),.o(intermediate_reg_1[2407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4813]),.i2(intermediate_reg_0[4812]),.o(intermediate_reg_1[2406])); 
fsm fsm_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4811]),.i2(intermediate_reg_0[4810]),.o(intermediate_reg_1[2405])); 
fsm fsm_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4809]),.i2(intermediate_reg_0[4808]),.o(intermediate_reg_1[2404])); 
mux_module mux_module_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4807]),.i2(intermediate_reg_0[4806]),.o(intermediate_reg_1[2403]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4805]),.i2(intermediate_reg_0[4804]),.o(intermediate_reg_1[2402])); 
mux_module mux_module_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4803]),.i2(intermediate_reg_0[4802]),.o(intermediate_reg_1[2401]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4801]),.i2(intermediate_reg_0[4800]),.o(intermediate_reg_1[2400]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4799]),.i2(intermediate_reg_0[4798]),.o(intermediate_reg_1[2399]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4797]),.i2(intermediate_reg_0[4796]),.o(intermediate_reg_1[2398])); 
mux_module mux_module_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4795]),.i2(intermediate_reg_0[4794]),.o(intermediate_reg_1[2397]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4793]),.i2(intermediate_reg_0[4792]),.o(intermediate_reg_1[2396])); 
mux_module mux_module_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4791]),.i2(intermediate_reg_0[4790]),.o(intermediate_reg_1[2395]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4789]),.i2(intermediate_reg_0[4788]),.o(intermediate_reg_1[2394]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4787]),.i2(intermediate_reg_0[4786]),.o(intermediate_reg_1[2393])); 
fsm fsm_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4785]),.i2(intermediate_reg_0[4784]),.o(intermediate_reg_1[2392])); 
mux_module mux_module_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4783]),.i2(intermediate_reg_0[4782]),.o(intermediate_reg_1[2391]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4781]),.i2(intermediate_reg_0[4780]),.o(intermediate_reg_1[2390]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4779]),.i2(intermediate_reg_0[4778]),.o(intermediate_reg_1[2389])); 
mux_module mux_module_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4777]),.i2(intermediate_reg_0[4776]),.o(intermediate_reg_1[2388]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4775]),.i2(intermediate_reg_0[4774]),.o(intermediate_reg_1[2387]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4773]),.i2(intermediate_reg_0[4772]),.o(intermediate_reg_1[2386])); 
mux_module mux_module_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4771]),.i2(intermediate_reg_0[4770]),.o(intermediate_reg_1[2385]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4769]),.i2(intermediate_reg_0[4768]),.o(intermediate_reg_1[2384])); 
mux_module mux_module_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4767]),.i2(intermediate_reg_0[4766]),.o(intermediate_reg_1[2383]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4765]),.i2(intermediate_reg_0[4764]),.o(intermediate_reg_1[2382])); 
fsm fsm_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4763]),.i2(intermediate_reg_0[4762]),.o(intermediate_reg_1[2381])); 
fsm fsm_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4761]),.i2(intermediate_reg_0[4760]),.o(intermediate_reg_1[2380])); 
mux_module mux_module_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4759]),.i2(intermediate_reg_0[4758]),.o(intermediate_reg_1[2379]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4757]),.i2(intermediate_reg_0[4756]),.o(intermediate_reg_1[2378])); 
mux_module mux_module_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4755]),.i2(intermediate_reg_0[4754]),.o(intermediate_reg_1[2377]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4753]),.i2(intermediate_reg_0[4752]),.o(intermediate_reg_1[2376])); 
fsm fsm_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4751]),.i2(intermediate_reg_0[4750]),.o(intermediate_reg_1[2375])); 
mux_module mux_module_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4749]),.i2(intermediate_reg_0[4748]),.o(intermediate_reg_1[2374]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4747]),.i2(intermediate_reg_0[4746]),.o(intermediate_reg_1[2373]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4745]),.i2(intermediate_reg_0[4744]),.o(intermediate_reg_1[2372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4743]),.i2(intermediate_reg_0[4742]),.o(intermediate_reg_1[2371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4741]),.i2(intermediate_reg_0[4740]),.o(intermediate_reg_1[2370]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4739]),.i2(intermediate_reg_0[4738]),.o(intermediate_reg_1[2369])); 
mux_module mux_module_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4737]),.i2(intermediate_reg_0[4736]),.o(intermediate_reg_1[2368]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4735]),.i2(intermediate_reg_0[4734]),.o(intermediate_reg_1[2367])); 
fsm fsm_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4733]),.i2(intermediate_reg_0[4732]),.o(intermediate_reg_1[2366])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4731]),.i2(intermediate_reg_0[4730]),.o(intermediate_reg_1[2365]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4729]),.i2(intermediate_reg_0[4728]),.o(intermediate_reg_1[2364])); 
mux_module mux_module_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4727]),.i2(intermediate_reg_0[4726]),.o(intermediate_reg_1[2363]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4725]),.i2(intermediate_reg_0[4724]),.o(intermediate_reg_1[2362]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4723]),.i2(intermediate_reg_0[4722]),.o(intermediate_reg_1[2361])); 
fsm fsm_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4721]),.i2(intermediate_reg_0[4720]),.o(intermediate_reg_1[2360])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4719]),.i2(intermediate_reg_0[4718]),.o(intermediate_reg_1[2359]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4717]),.i2(intermediate_reg_0[4716]),.o(intermediate_reg_1[2358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4715]),.i2(intermediate_reg_0[4714]),.o(intermediate_reg_1[2357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4713]),.i2(intermediate_reg_0[4712]),.o(intermediate_reg_1[2356]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4711]),.i2(intermediate_reg_0[4710]),.o(intermediate_reg_1[2355])); 
mux_module mux_module_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4709]),.i2(intermediate_reg_0[4708]),.o(intermediate_reg_1[2354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4707]),.i2(intermediate_reg_0[4706]),.o(intermediate_reg_1[2353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4705]),.i2(intermediate_reg_0[4704]),.o(intermediate_reg_1[2352]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4703]),.i2(intermediate_reg_0[4702]),.o(intermediate_reg_1[2351])); 
fsm fsm_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4701]),.i2(intermediate_reg_0[4700]),.o(intermediate_reg_1[2350])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4699]),.i2(intermediate_reg_0[4698]),.o(intermediate_reg_1[2349]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4697]),.i2(intermediate_reg_0[4696]),.o(intermediate_reg_1[2348]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4695]),.i2(intermediate_reg_0[4694]),.o(intermediate_reg_1[2347])); 
mux_module mux_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4693]),.i2(intermediate_reg_0[4692]),.o(intermediate_reg_1[2346]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4691]),.i2(intermediate_reg_0[4690]),.o(intermediate_reg_1[2345]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4689]),.i2(intermediate_reg_0[4688]),.o(intermediate_reg_1[2344])); 
fsm fsm_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4687]),.i2(intermediate_reg_0[4686]),.o(intermediate_reg_1[2343])); 
fsm fsm_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4685]),.i2(intermediate_reg_0[4684]),.o(intermediate_reg_1[2342])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4683]),.i2(intermediate_reg_0[4682]),.o(intermediate_reg_1[2341]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4681]),.i2(intermediate_reg_0[4680]),.o(intermediate_reg_1[2340]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4679]),.i2(intermediate_reg_0[4678]),.o(intermediate_reg_1[2339]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4677]),.i2(intermediate_reg_0[4676]),.o(intermediate_reg_1[2338])); 
mux_module mux_module_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4675]),.i2(intermediate_reg_0[4674]),.o(intermediate_reg_1[2337]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4673]),.i2(intermediate_reg_0[4672]),.o(intermediate_reg_1[2336])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4671]),.i2(intermediate_reg_0[4670]),.o(intermediate_reg_1[2335])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4669]),.i2(intermediate_reg_0[4668]),.o(intermediate_reg_1[2334])); 
fsm fsm_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4667]),.i2(intermediate_reg_0[4666]),.o(intermediate_reg_1[2333])); 
fsm fsm_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4665]),.i2(intermediate_reg_0[4664]),.o(intermediate_reg_1[2332])); 
mux_module mux_module_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4663]),.i2(intermediate_reg_0[4662]),.o(intermediate_reg_1[2331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4661]),.i2(intermediate_reg_0[4660]),.o(intermediate_reg_1[2330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4659]),.i2(intermediate_reg_0[4658]),.o(intermediate_reg_1[2329]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4657]),.i2(intermediate_reg_0[4656]),.o(intermediate_reg_1[2328])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4655]),.i2(intermediate_reg_0[4654]),.o(intermediate_reg_1[2327]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4653]),.i2(intermediate_reg_0[4652]),.o(intermediate_reg_1[2326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4651]),.i2(intermediate_reg_0[4650]),.o(intermediate_reg_1[2325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4649]),.i2(intermediate_reg_0[4648]),.o(intermediate_reg_1[2324]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4647]),.i2(intermediate_reg_0[4646]),.o(intermediate_reg_1[2323])); 
fsm fsm_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4645]),.i2(intermediate_reg_0[4644]),.o(intermediate_reg_1[2322])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4643]),.i2(intermediate_reg_0[4642]),.o(intermediate_reg_1[2321])); 
fsm fsm_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4641]),.i2(intermediate_reg_0[4640]),.o(intermediate_reg_1[2320])); 
mux_module mux_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4639]),.i2(intermediate_reg_0[4638]),.o(intermediate_reg_1[2319]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4637]),.i2(intermediate_reg_0[4636]),.o(intermediate_reg_1[2318])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4635]),.i2(intermediate_reg_0[4634]),.o(intermediate_reg_1[2317])); 
fsm fsm_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4633]),.i2(intermediate_reg_0[4632]),.o(intermediate_reg_1[2316])); 
fsm fsm_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4631]),.i2(intermediate_reg_0[4630]),.o(intermediate_reg_1[2315])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4629]),.i2(intermediate_reg_0[4628]),.o(intermediate_reg_1[2314]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4627]),.i2(intermediate_reg_0[4626]),.o(intermediate_reg_1[2313]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4625]),.i2(intermediate_reg_0[4624]),.o(intermediate_reg_1[2312])); 
mux_module mux_module_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4623]),.i2(intermediate_reg_0[4622]),.o(intermediate_reg_1[2311]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4621]),.i2(intermediate_reg_0[4620]),.o(intermediate_reg_1[2310]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4619]),.i2(intermediate_reg_0[4618]),.o(intermediate_reg_1[2309])); 
fsm fsm_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4617]),.i2(intermediate_reg_0[4616]),.o(intermediate_reg_1[2308])); 
fsm fsm_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4615]),.i2(intermediate_reg_0[4614]),.o(intermediate_reg_1[2307])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4613]),.i2(intermediate_reg_0[4612]),.o(intermediate_reg_1[2306]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4611]),.i2(intermediate_reg_0[4610]),.o(intermediate_reg_1[2305])); 
mux_module mux_module_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4609]),.i2(intermediate_reg_0[4608]),.o(intermediate_reg_1[2304]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4607]),.i2(intermediate_reg_0[4606]),.o(intermediate_reg_1[2303])); 
fsm fsm_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4605]),.i2(intermediate_reg_0[4604]),.o(intermediate_reg_1[2302])); 
mux_module mux_module_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4603]),.i2(intermediate_reg_0[4602]),.o(intermediate_reg_1[2301]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4601]),.i2(intermediate_reg_0[4600]),.o(intermediate_reg_1[2300])); 
mux_module mux_module_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4599]),.i2(intermediate_reg_0[4598]),.o(intermediate_reg_1[2299]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4597]),.i2(intermediate_reg_0[4596]),.o(intermediate_reg_1[2298])); 
fsm fsm_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4595]),.i2(intermediate_reg_0[4594]),.o(intermediate_reg_1[2297])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4593]),.i2(intermediate_reg_0[4592]),.o(intermediate_reg_1[2296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4591]),.i2(intermediate_reg_0[4590]),.o(intermediate_reg_1[2295]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4589]),.i2(intermediate_reg_0[4588]),.o(intermediate_reg_1[2294])); 
fsm fsm_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4587]),.i2(intermediate_reg_0[4586]),.o(intermediate_reg_1[2293])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4585]),.i2(intermediate_reg_0[4584]),.o(intermediate_reg_1[2292]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4583]),.i2(intermediate_reg_0[4582]),.o(intermediate_reg_1[2291])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4581]),.i2(intermediate_reg_0[4580]),.o(intermediate_reg_1[2290]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4579]),.i2(intermediate_reg_0[4578]),.o(intermediate_reg_1[2289]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4577]),.i2(intermediate_reg_0[4576]),.o(intermediate_reg_1[2288]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4575]),.i2(intermediate_reg_0[4574]),.o(intermediate_reg_1[2287])); 
fsm fsm_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4573]),.i2(intermediate_reg_0[4572]),.o(intermediate_reg_1[2286])); 
fsm fsm_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4571]),.i2(intermediate_reg_0[4570]),.o(intermediate_reg_1[2285])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4569]),.i2(intermediate_reg_0[4568]),.o(intermediate_reg_1[2284]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4567]),.i2(intermediate_reg_0[4566]),.o(intermediate_reg_1[2283])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4565]),.i2(intermediate_reg_0[4564]),.o(intermediate_reg_1[2282])); 
fsm fsm_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4563]),.i2(intermediate_reg_0[4562]),.o(intermediate_reg_1[2281])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4561]),.i2(intermediate_reg_0[4560]),.o(intermediate_reg_1[2280])); 
mux_module mux_module_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4559]),.i2(intermediate_reg_0[4558]),.o(intermediate_reg_1[2279]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4557]),.i2(intermediate_reg_0[4556]),.o(intermediate_reg_1[2278]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4555]),.i2(intermediate_reg_0[4554]),.o(intermediate_reg_1[2277]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4553]),.i2(intermediate_reg_0[4552]),.o(intermediate_reg_1[2276])); 
fsm fsm_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4551]),.i2(intermediate_reg_0[4550]),.o(intermediate_reg_1[2275])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4549]),.i2(intermediate_reg_0[4548]),.o(intermediate_reg_1[2274])); 
fsm fsm_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4547]),.i2(intermediate_reg_0[4546]),.o(intermediate_reg_1[2273])); 
mux_module mux_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4545]),.i2(intermediate_reg_0[4544]),.o(intermediate_reg_1[2272]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4543]),.i2(intermediate_reg_0[4542]),.o(intermediate_reg_1[2271])); 
fsm fsm_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4541]),.i2(intermediate_reg_0[4540]),.o(intermediate_reg_1[2270])); 
fsm fsm_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4539]),.i2(intermediate_reg_0[4538]),.o(intermediate_reg_1[2269])); 
mux_module mux_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4537]),.i2(intermediate_reg_0[4536]),.o(intermediate_reg_1[2268]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4535]),.i2(intermediate_reg_0[4534]),.o(intermediate_reg_1[2267]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4533]),.i2(intermediate_reg_0[4532]),.o(intermediate_reg_1[2266])); 
fsm fsm_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4531]),.i2(intermediate_reg_0[4530]),.o(intermediate_reg_1[2265])); 
mux_module mux_module_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4529]),.i2(intermediate_reg_0[4528]),.o(intermediate_reg_1[2264]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4527]),.i2(intermediate_reg_0[4526]),.o(intermediate_reg_1[2263]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4525]),.i2(intermediate_reg_0[4524]),.o(intermediate_reg_1[2262])); 
fsm fsm_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4523]),.i2(intermediate_reg_0[4522]),.o(intermediate_reg_1[2261])); 
fsm fsm_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4521]),.i2(intermediate_reg_0[4520]),.o(intermediate_reg_1[2260])); 
fsm fsm_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4519]),.i2(intermediate_reg_0[4518]),.o(intermediate_reg_1[2259])); 
fsm fsm_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4517]),.i2(intermediate_reg_0[4516]),.o(intermediate_reg_1[2258])); 
fsm fsm_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4515]),.i2(intermediate_reg_0[4514]),.o(intermediate_reg_1[2257])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4513]),.i2(intermediate_reg_0[4512]),.o(intermediate_reg_1[2256])); 
mux_module mux_module_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4511]),.i2(intermediate_reg_0[4510]),.o(intermediate_reg_1[2255]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4509]),.i2(intermediate_reg_0[4508]),.o(intermediate_reg_1[2254])); 
mux_module mux_module_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4507]),.i2(intermediate_reg_0[4506]),.o(intermediate_reg_1[2253]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4505]),.i2(intermediate_reg_0[4504]),.o(intermediate_reg_1[2252])); 
mux_module mux_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4503]),.i2(intermediate_reg_0[4502]),.o(intermediate_reg_1[2251]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4501]),.i2(intermediate_reg_0[4500]),.o(intermediate_reg_1[2250])); 
mux_module mux_module_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4499]),.i2(intermediate_reg_0[4498]),.o(intermediate_reg_1[2249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4497]),.i2(intermediate_reg_0[4496]),.o(intermediate_reg_1[2248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4495]),.i2(intermediate_reg_0[4494]),.o(intermediate_reg_1[2247]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4493]),.i2(intermediate_reg_0[4492]),.o(intermediate_reg_1[2246])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4491]),.i2(intermediate_reg_0[4490]),.o(intermediate_reg_1[2245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4489]),.i2(intermediate_reg_0[4488]),.o(intermediate_reg_1[2244]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4487]),.i2(intermediate_reg_0[4486]),.o(intermediate_reg_1[2243]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4485]),.i2(intermediate_reg_0[4484]),.o(intermediate_reg_1[2242])); 
fsm fsm_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4483]),.i2(intermediate_reg_0[4482]),.o(intermediate_reg_1[2241])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4481]),.i2(intermediate_reg_0[4480]),.o(intermediate_reg_1[2240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4479]),.i2(intermediate_reg_0[4478]),.o(intermediate_reg_1[2239]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4477]),.i2(intermediate_reg_0[4476]),.o(intermediate_reg_1[2238])); 
fsm fsm_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4475]),.i2(intermediate_reg_0[4474]),.o(intermediate_reg_1[2237])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4473]),.i2(intermediate_reg_0[4472]),.o(intermediate_reg_1[2236]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4471]),.i2(intermediate_reg_0[4470]),.o(intermediate_reg_1[2235])); 
mux_module mux_module_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4469]),.i2(intermediate_reg_0[4468]),.o(intermediate_reg_1[2234]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4467]),.i2(intermediate_reg_0[4466]),.o(intermediate_reg_1[2233])); 
fsm fsm_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4465]),.i2(intermediate_reg_0[4464]),.o(intermediate_reg_1[2232])); 
fsm fsm_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4463]),.i2(intermediate_reg_0[4462]),.o(intermediate_reg_1[2231])); 
mux_module mux_module_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4461]),.i2(intermediate_reg_0[4460]),.o(intermediate_reg_1[2230]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4459]),.i2(intermediate_reg_0[4458]),.o(intermediate_reg_1[2229])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4457]),.i2(intermediate_reg_0[4456]),.o(intermediate_reg_1[2228])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4455]),.i2(intermediate_reg_0[4454]),.o(intermediate_reg_1[2227]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4453]),.i2(intermediate_reg_0[4452]),.o(intermediate_reg_1[2226])); 
fsm fsm_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4451]),.i2(intermediate_reg_0[4450]),.o(intermediate_reg_1[2225])); 
mux_module mux_module_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4449]),.i2(intermediate_reg_0[4448]),.o(intermediate_reg_1[2224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4447]),.i2(intermediate_reg_0[4446]),.o(intermediate_reg_1[2223]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4445]),.i2(intermediate_reg_0[4444]),.o(intermediate_reg_1[2222])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4443]),.i2(intermediate_reg_0[4442]),.o(intermediate_reg_1[2221])); 
fsm fsm_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4441]),.i2(intermediate_reg_0[4440]),.o(intermediate_reg_1[2220])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4439]),.i2(intermediate_reg_0[4438]),.o(intermediate_reg_1[2219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4437]),.i2(intermediate_reg_0[4436]),.o(intermediate_reg_1[2218]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4435]),.i2(intermediate_reg_0[4434]),.o(intermediate_reg_1[2217])); 
fsm fsm_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4433]),.i2(intermediate_reg_0[4432]),.o(intermediate_reg_1[2216])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4431]),.i2(intermediate_reg_0[4430]),.o(intermediate_reg_1[2215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4429]),.i2(intermediate_reg_0[4428]),.o(intermediate_reg_1[2214]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4427]),.i2(intermediate_reg_0[4426]),.o(intermediate_reg_1[2213])); 
mux_module mux_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4425]),.i2(intermediate_reg_0[4424]),.o(intermediate_reg_1[2212]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4423]),.i2(intermediate_reg_0[4422]),.o(intermediate_reg_1[2211]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4421]),.i2(intermediate_reg_0[4420]),.o(intermediate_reg_1[2210]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4419]),.i2(intermediate_reg_0[4418]),.o(intermediate_reg_1[2209])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4417]),.i2(intermediate_reg_0[4416]),.o(intermediate_reg_1[2208]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4415]),.i2(intermediate_reg_0[4414]),.o(intermediate_reg_1[2207])); 
mux_module mux_module_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4413]),.i2(intermediate_reg_0[4412]),.o(intermediate_reg_1[2206]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4411]),.i2(intermediate_reg_0[4410]),.o(intermediate_reg_1[2205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4409]),.i2(intermediate_reg_0[4408]),.o(intermediate_reg_1[2204]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4407]),.i2(intermediate_reg_0[4406]),.o(intermediate_reg_1[2203])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4405]),.i2(intermediate_reg_0[4404]),.o(intermediate_reg_1[2202])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4403]),.i2(intermediate_reg_0[4402]),.o(intermediate_reg_1[2201]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4401]),.i2(intermediate_reg_0[4400]),.o(intermediate_reg_1[2200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4399]),.i2(intermediate_reg_0[4398]),.o(intermediate_reg_1[2199]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4397]),.i2(intermediate_reg_0[4396]),.o(intermediate_reg_1[2198]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4395]),.i2(intermediate_reg_0[4394]),.o(intermediate_reg_1[2197])); 
mux_module mux_module_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4393]),.i2(intermediate_reg_0[4392]),.o(intermediate_reg_1[2196]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4391]),.i2(intermediate_reg_0[4390]),.o(intermediate_reg_1[2195])); 
mux_module mux_module_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4389]),.i2(intermediate_reg_0[4388]),.o(intermediate_reg_1[2194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4387]),.i2(intermediate_reg_0[4386]),.o(intermediate_reg_1[2193]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4385]),.i2(intermediate_reg_0[4384]),.o(intermediate_reg_1[2192])); 
mux_module mux_module_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4383]),.i2(intermediate_reg_0[4382]),.o(intermediate_reg_1[2191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4381]),.i2(intermediate_reg_0[4380]),.o(intermediate_reg_1[2190]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4379]),.i2(intermediate_reg_0[4378]),.o(intermediate_reg_1[2189])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4377]),.i2(intermediate_reg_0[4376]),.o(intermediate_reg_1[2188])); 
mux_module mux_module_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4375]),.i2(intermediate_reg_0[4374]),.o(intermediate_reg_1[2187]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4373]),.i2(intermediate_reg_0[4372]),.o(intermediate_reg_1[2186]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4371]),.i2(intermediate_reg_0[4370]),.o(intermediate_reg_1[2185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4369]),.i2(intermediate_reg_0[4368]),.o(intermediate_reg_1[2184]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4367]),.i2(intermediate_reg_0[4366]),.o(intermediate_reg_1[2183]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4365]),.i2(intermediate_reg_0[4364]),.o(intermediate_reg_1[2182]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4363]),.i2(intermediate_reg_0[4362]),.o(intermediate_reg_1[2181])); 
mux_module mux_module_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4361]),.i2(intermediate_reg_0[4360]),.o(intermediate_reg_1[2180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4359]),.i2(intermediate_reg_0[4358]),.o(intermediate_reg_1[2179]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4357]),.i2(intermediate_reg_0[4356]),.o(intermediate_reg_1[2178])); 
fsm fsm_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4355]),.i2(intermediate_reg_0[4354]),.o(intermediate_reg_1[2177])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4353]),.i2(intermediate_reg_0[4352]),.o(intermediate_reg_1[2176])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4351]),.i2(intermediate_reg_0[4350]),.o(intermediate_reg_1[2175])); 
fsm fsm_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4349]),.i2(intermediate_reg_0[4348]),.o(intermediate_reg_1[2174])); 
mux_module mux_module_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4347]),.i2(intermediate_reg_0[4346]),.o(intermediate_reg_1[2173]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4345]),.i2(intermediate_reg_0[4344]),.o(intermediate_reg_1[2172])); 
fsm fsm_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4343]),.i2(intermediate_reg_0[4342]),.o(intermediate_reg_1[2171])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4341]),.i2(intermediate_reg_0[4340]),.o(intermediate_reg_1[2170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4339]),.i2(intermediate_reg_0[4338]),.o(intermediate_reg_1[2169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4337]),.i2(intermediate_reg_0[4336]),.o(intermediate_reg_1[2168]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4335]),.i2(intermediate_reg_0[4334]),.o(intermediate_reg_1[2167]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4333]),.i2(intermediate_reg_0[4332]),.o(intermediate_reg_1[2166]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4331]),.i2(intermediate_reg_0[4330]),.o(intermediate_reg_1[2165]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4329]),.i2(intermediate_reg_0[4328]),.o(intermediate_reg_1[2164]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4327]),.i2(intermediate_reg_0[4326]),.o(intermediate_reg_1[2163])); 
fsm fsm_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4325]),.i2(intermediate_reg_0[4324]),.o(intermediate_reg_1[2162])); 
mux_module mux_module_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4323]),.i2(intermediate_reg_0[4322]),.o(intermediate_reg_1[2161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4321]),.i2(intermediate_reg_0[4320]),.o(intermediate_reg_1[2160]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4319]),.i2(intermediate_reg_0[4318]),.o(intermediate_reg_1[2159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4317]),.i2(intermediate_reg_0[4316]),.o(intermediate_reg_1[2158]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4315]),.i2(intermediate_reg_0[4314]),.o(intermediate_reg_1[2157])); 
fsm fsm_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4313]),.i2(intermediate_reg_0[4312]),.o(intermediate_reg_1[2156])); 
fsm fsm_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4311]),.i2(intermediate_reg_0[4310]),.o(intermediate_reg_1[2155])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4309]),.i2(intermediate_reg_0[4308]),.o(intermediate_reg_1[2154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4307]),.i2(intermediate_reg_0[4306]),.o(intermediate_reg_1[2153]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4305]),.i2(intermediate_reg_0[4304]),.o(intermediate_reg_1[2152])); 
fsm fsm_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4303]),.i2(intermediate_reg_0[4302]),.o(intermediate_reg_1[2151])); 
mux_module mux_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4301]),.i2(intermediate_reg_0[4300]),.o(intermediate_reg_1[2150]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4299]),.i2(intermediate_reg_0[4298]),.o(intermediate_reg_1[2149]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4297]),.i2(intermediate_reg_0[4296]),.o(intermediate_reg_1[2148])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4295]),.i2(intermediate_reg_0[4294]),.o(intermediate_reg_1[2147]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4293]),.i2(intermediate_reg_0[4292]),.o(intermediate_reg_1[2146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4291]),.i2(intermediate_reg_0[4290]),.o(intermediate_reg_1[2145]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4289]),.i2(intermediate_reg_0[4288]),.o(intermediate_reg_1[2144])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4287]),.i2(intermediate_reg_0[4286]),.o(intermediate_reg_1[2143]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4285]),.i2(intermediate_reg_0[4284]),.o(intermediate_reg_1[2142]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4283]),.i2(intermediate_reg_0[4282]),.o(intermediate_reg_1[2141])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4281]),.i2(intermediate_reg_0[4280]),.o(intermediate_reg_1[2140]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4279]),.i2(intermediate_reg_0[4278]),.o(intermediate_reg_1[2139]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4277]),.i2(intermediate_reg_0[4276]),.o(intermediate_reg_1[2138])); 
fsm fsm_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4275]),.i2(intermediate_reg_0[4274]),.o(intermediate_reg_1[2137])); 
fsm fsm_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4273]),.i2(intermediate_reg_0[4272]),.o(intermediate_reg_1[2136])); 
mux_module mux_module_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4271]),.i2(intermediate_reg_0[4270]),.o(intermediate_reg_1[2135]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4269]),.i2(intermediate_reg_0[4268]),.o(intermediate_reg_1[2134])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4267]),.i2(intermediate_reg_0[4266]),.o(intermediate_reg_1[2133])); 
mux_module mux_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4265]),.i2(intermediate_reg_0[4264]),.o(intermediate_reg_1[2132]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4263]),.i2(intermediate_reg_0[4262]),.o(intermediate_reg_1[2131])); 
mux_module mux_module_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4261]),.i2(intermediate_reg_0[4260]),.o(intermediate_reg_1[2130]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4259]),.i2(intermediate_reg_0[4258]),.o(intermediate_reg_1[2129]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4257]),.i2(intermediate_reg_0[4256]),.o(intermediate_reg_1[2128]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4255]),.i2(intermediate_reg_0[4254]),.o(intermediate_reg_1[2127])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4253]),.i2(intermediate_reg_0[4252]),.o(intermediate_reg_1[2126])); 
fsm fsm_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4251]),.i2(intermediate_reg_0[4250]),.o(intermediate_reg_1[2125])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4249]),.i2(intermediate_reg_0[4248]),.o(intermediate_reg_1[2124]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4247]),.i2(intermediate_reg_0[4246]),.o(intermediate_reg_1[2123]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4245]),.i2(intermediate_reg_0[4244]),.o(intermediate_reg_1[2122]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4243]),.i2(intermediate_reg_0[4242]),.o(intermediate_reg_1[2121])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4241]),.i2(intermediate_reg_0[4240]),.o(intermediate_reg_1[2120])); 
fsm fsm_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4239]),.i2(intermediate_reg_0[4238]),.o(intermediate_reg_1[2119])); 
mux_module mux_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4237]),.i2(intermediate_reg_0[4236]),.o(intermediate_reg_1[2118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4235]),.i2(intermediate_reg_0[4234]),.o(intermediate_reg_1[2117]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4233]),.i2(intermediate_reg_0[4232]),.o(intermediate_reg_1[2116])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4231]),.i2(intermediate_reg_0[4230]),.o(intermediate_reg_1[2115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4229]),.i2(intermediate_reg_0[4228]),.o(intermediate_reg_1[2114])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4227]),.i2(intermediate_reg_0[4226]),.o(intermediate_reg_1[2113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4225]),.i2(intermediate_reg_0[4224]),.o(intermediate_reg_1[2112]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4223]),.i2(intermediate_reg_0[4222]),.o(intermediate_reg_1[2111])); 
fsm fsm_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4221]),.i2(intermediate_reg_0[4220]),.o(intermediate_reg_1[2110])); 
fsm fsm_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4219]),.i2(intermediate_reg_0[4218]),.o(intermediate_reg_1[2109])); 
fsm fsm_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4217]),.i2(intermediate_reg_0[4216]),.o(intermediate_reg_1[2108])); 
fsm fsm_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4215]),.i2(intermediate_reg_0[4214]),.o(intermediate_reg_1[2107])); 
mux_module mux_module_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4213]),.i2(intermediate_reg_0[4212]),.o(intermediate_reg_1[2106]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4211]),.i2(intermediate_reg_0[4210]),.o(intermediate_reg_1[2105])); 
fsm fsm_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4209]),.i2(intermediate_reg_0[4208]),.o(intermediate_reg_1[2104])); 
mux_module mux_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4207]),.i2(intermediate_reg_0[4206]),.o(intermediate_reg_1[2103]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4205]),.i2(intermediate_reg_0[4204]),.o(intermediate_reg_1[2102])); 
fsm fsm_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4203]),.i2(intermediate_reg_0[4202]),.o(intermediate_reg_1[2101])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4201]),.i2(intermediate_reg_0[4200]),.o(intermediate_reg_1[2100])); 
mux_module mux_module_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4199]),.i2(intermediate_reg_0[4198]),.o(intermediate_reg_1[2099]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4197]),.i2(intermediate_reg_0[4196]),.o(intermediate_reg_1[2098])); 
mux_module mux_module_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4195]),.i2(intermediate_reg_0[4194]),.o(intermediate_reg_1[2097]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4193]),.i2(intermediate_reg_0[4192]),.o(intermediate_reg_1[2096])); 
fsm fsm_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4191]),.i2(intermediate_reg_0[4190]),.o(intermediate_reg_1[2095])); 
mux_module mux_module_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4189]),.i2(intermediate_reg_0[4188]),.o(intermediate_reg_1[2094]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4187]),.i2(intermediate_reg_0[4186]),.o(intermediate_reg_1[2093])); 
mux_module mux_module_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4185]),.i2(intermediate_reg_0[4184]),.o(intermediate_reg_1[2092]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4183]),.i2(intermediate_reg_0[4182]),.o(intermediate_reg_1[2091]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4181]),.i2(intermediate_reg_0[4180]),.o(intermediate_reg_1[2090]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4179]),.i2(intermediate_reg_0[4178]),.o(intermediate_reg_1[2089])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4177]),.i2(intermediate_reg_0[4176]),.o(intermediate_reg_1[2088])); 
mux_module mux_module_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4175]),.i2(intermediate_reg_0[4174]),.o(intermediate_reg_1[2087]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4173]),.i2(intermediate_reg_0[4172]),.o(intermediate_reg_1[2086]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4171]),.i2(intermediate_reg_0[4170]),.o(intermediate_reg_1[2085])); 
fsm fsm_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4169]),.i2(intermediate_reg_0[4168]),.o(intermediate_reg_1[2084])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4167]),.i2(intermediate_reg_0[4166]),.o(intermediate_reg_1[2083]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4165]),.i2(intermediate_reg_0[4164]),.o(intermediate_reg_1[2082])); 
fsm fsm_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4163]),.i2(intermediate_reg_0[4162]),.o(intermediate_reg_1[2081])); 
fsm fsm_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4161]),.i2(intermediate_reg_0[4160]),.o(intermediate_reg_1[2080])); 
mux_module mux_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4159]),.i2(intermediate_reg_0[4158]),.o(intermediate_reg_1[2079]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4157]),.i2(intermediate_reg_0[4156]),.o(intermediate_reg_1[2078]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4155]),.i2(intermediate_reg_0[4154]),.o(intermediate_reg_1[2077]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4153]),.i2(intermediate_reg_0[4152]),.o(intermediate_reg_1[2076]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4151]),.i2(intermediate_reg_0[4150]),.o(intermediate_reg_1[2075])); 
fsm fsm_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4149]),.i2(intermediate_reg_0[4148]),.o(intermediate_reg_1[2074])); 
mux_module mux_module_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4147]),.i2(intermediate_reg_0[4146]),.o(intermediate_reg_1[2073]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4145]),.i2(intermediate_reg_0[4144]),.o(intermediate_reg_1[2072]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4143]),.i2(intermediate_reg_0[4142]),.o(intermediate_reg_1[2071])); 
fsm fsm_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4141]),.i2(intermediate_reg_0[4140]),.o(intermediate_reg_1[2070])); 
fsm fsm_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4139]),.i2(intermediate_reg_0[4138]),.o(intermediate_reg_1[2069])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4137]),.i2(intermediate_reg_0[4136]),.o(intermediate_reg_1[2068]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4135]),.i2(intermediate_reg_0[4134]),.o(intermediate_reg_1[2067]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4133]),.i2(intermediate_reg_0[4132]),.o(intermediate_reg_1[2066])); 
fsm fsm_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4131]),.i2(intermediate_reg_0[4130]),.o(intermediate_reg_1[2065])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4129]),.i2(intermediate_reg_0[4128]),.o(intermediate_reg_1[2064]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4127]),.i2(intermediate_reg_0[4126]),.o(intermediate_reg_1[2063])); 
fsm fsm_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4125]),.i2(intermediate_reg_0[4124]),.o(intermediate_reg_1[2062])); 
mux_module mux_module_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4123]),.i2(intermediate_reg_0[4122]),.o(intermediate_reg_1[2061]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4121]),.i2(intermediate_reg_0[4120]),.o(intermediate_reg_1[2060])); 
fsm fsm_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4119]),.i2(intermediate_reg_0[4118]),.o(intermediate_reg_1[2059])); 
fsm fsm_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4117]),.i2(intermediate_reg_0[4116]),.o(intermediate_reg_1[2058])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4115]),.i2(intermediate_reg_0[4114]),.o(intermediate_reg_1[2057]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4113]),.i2(intermediate_reg_0[4112]),.o(intermediate_reg_1[2056]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4111]),.i2(intermediate_reg_0[4110]),.o(intermediate_reg_1[2055]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4109]),.i2(intermediate_reg_0[4108]),.o(intermediate_reg_1[2054]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4107]),.i2(intermediate_reg_0[4106]),.o(intermediate_reg_1[2053]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4105]),.i2(intermediate_reg_0[4104]),.o(intermediate_reg_1[2052])); 
mux_module mux_module_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4103]),.i2(intermediate_reg_0[4102]),.o(intermediate_reg_1[2051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4101]),.i2(intermediate_reg_0[4100]),.o(intermediate_reg_1[2050]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4099]),.i2(intermediate_reg_0[4098]),.o(intermediate_reg_1[2049]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4097]),.i2(intermediate_reg_0[4096]),.o(intermediate_reg_1[2048]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4095]),.i2(intermediate_reg_0[4094]),.o(intermediate_reg_1[2047])); 
fsm fsm_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4093]),.i2(intermediate_reg_0[4092]),.o(intermediate_reg_1[2046])); 
fsm fsm_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4091]),.i2(intermediate_reg_0[4090]),.o(intermediate_reg_1[2045])); 
mux_module mux_module_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4089]),.i2(intermediate_reg_0[4088]),.o(intermediate_reg_1[2044]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4087]),.i2(intermediate_reg_0[4086]),.o(intermediate_reg_1[2043]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4085]),.i2(intermediate_reg_0[4084]),.o(intermediate_reg_1[2042]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4083]),.i2(intermediate_reg_0[4082]),.o(intermediate_reg_1[2041]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4081]),.i2(intermediate_reg_0[4080]),.o(intermediate_reg_1[2040])); 
fsm fsm_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4079]),.i2(intermediate_reg_0[4078]),.o(intermediate_reg_1[2039])); 
fsm fsm_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4077]),.i2(intermediate_reg_0[4076]),.o(intermediate_reg_1[2038])); 
mux_module mux_module_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4075]),.i2(intermediate_reg_0[4074]),.o(intermediate_reg_1[2037]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4073]),.i2(intermediate_reg_0[4072]),.o(intermediate_reg_1[2036])); 
fsm fsm_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4071]),.i2(intermediate_reg_0[4070]),.o(intermediate_reg_1[2035])); 
fsm fsm_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4069]),.i2(intermediate_reg_0[4068]),.o(intermediate_reg_1[2034])); 
fsm fsm_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4067]),.i2(intermediate_reg_0[4066]),.o(intermediate_reg_1[2033])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4065]),.i2(intermediate_reg_0[4064]),.o(intermediate_reg_1[2032]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4063]),.i2(intermediate_reg_0[4062]),.o(intermediate_reg_1[2031])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4061]),.i2(intermediate_reg_0[4060]),.o(intermediate_reg_1[2030]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4059]),.i2(intermediate_reg_0[4058]),.o(intermediate_reg_1[2029])); 
fsm fsm_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4057]),.i2(intermediate_reg_0[4056]),.o(intermediate_reg_1[2028])); 
mux_module mux_module_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4055]),.i2(intermediate_reg_0[4054]),.o(intermediate_reg_1[2027]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4053]),.i2(intermediate_reg_0[4052]),.o(intermediate_reg_1[2026]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4051]),.i2(intermediate_reg_0[4050]),.o(intermediate_reg_1[2025])); 
fsm fsm_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4049]),.i2(intermediate_reg_0[4048]),.o(intermediate_reg_1[2024])); 
fsm fsm_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4047]),.i2(intermediate_reg_0[4046]),.o(intermediate_reg_1[2023])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4045]),.i2(intermediate_reg_0[4044]),.o(intermediate_reg_1[2022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4043]),.i2(intermediate_reg_0[4042]),.o(intermediate_reg_1[2021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4041]),.i2(intermediate_reg_0[4040]),.o(intermediate_reg_1[2020]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4039]),.i2(intermediate_reg_0[4038]),.o(intermediate_reg_1[2019])); 
fsm fsm_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4037]),.i2(intermediate_reg_0[4036]),.o(intermediate_reg_1[2018])); 
fsm fsm_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4035]),.i2(intermediate_reg_0[4034]),.o(intermediate_reg_1[2017])); 
mux_module mux_module_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4033]),.i2(intermediate_reg_0[4032]),.o(intermediate_reg_1[2016]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4031]),.i2(intermediate_reg_0[4030]),.o(intermediate_reg_1[2015]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4029]),.i2(intermediate_reg_0[4028]),.o(intermediate_reg_1[2014])); 
fsm fsm_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4027]),.i2(intermediate_reg_0[4026]),.o(intermediate_reg_1[2013])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4025]),.i2(intermediate_reg_0[4024]),.o(intermediate_reg_1[2012])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4023]),.i2(intermediate_reg_0[4022]),.o(intermediate_reg_1[2011]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4021]),.i2(intermediate_reg_0[4020]),.o(intermediate_reg_1[2010])); 
fsm fsm_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4019]),.i2(intermediate_reg_0[4018]),.o(intermediate_reg_1[2009])); 
mux_module mux_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4017]),.i2(intermediate_reg_0[4016]),.o(intermediate_reg_1[2008]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4015]),.i2(intermediate_reg_0[4014]),.o(intermediate_reg_1[2007]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4013]),.i2(intermediate_reg_0[4012]),.o(intermediate_reg_1[2006])); 
fsm fsm_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4011]),.i2(intermediate_reg_0[4010]),.o(intermediate_reg_1[2005])); 
mux_module mux_module_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4009]),.i2(intermediate_reg_0[4008]),.o(intermediate_reg_1[2004]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4007]),.i2(intermediate_reg_0[4006]),.o(intermediate_reg_1[2003]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4005]),.i2(intermediate_reg_0[4004]),.o(intermediate_reg_1[2002])); 
mux_module mux_module_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4003]),.i2(intermediate_reg_0[4002]),.o(intermediate_reg_1[2001]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[4001]),.i2(intermediate_reg_0[4000]),.o(intermediate_reg_1[2000])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3999]),.i2(intermediate_reg_0[3998]),.o(intermediate_reg_1[1999]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3997]),.i2(intermediate_reg_0[3996]),.o(intermediate_reg_1[1998])); 
mux_module mux_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3995]),.i2(intermediate_reg_0[3994]),.o(intermediate_reg_1[1997]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3993]),.i2(intermediate_reg_0[3992]),.o(intermediate_reg_1[1996]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3991]),.i2(intermediate_reg_0[3990]),.o(intermediate_reg_1[1995])); 
fsm fsm_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3989]),.i2(intermediate_reg_0[3988]),.o(intermediate_reg_1[1994])); 
fsm fsm_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3987]),.i2(intermediate_reg_0[3986]),.o(intermediate_reg_1[1993])); 
mux_module mux_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3985]),.i2(intermediate_reg_0[3984]),.o(intermediate_reg_1[1992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3983]),.i2(intermediate_reg_0[3982]),.o(intermediate_reg_1[1991]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3981]),.i2(intermediate_reg_0[3980]),.o(intermediate_reg_1[1990])); 
mux_module mux_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3979]),.i2(intermediate_reg_0[3978]),.o(intermediate_reg_1[1989]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3977]),.i2(intermediate_reg_0[3976]),.o(intermediate_reg_1[1988])); 
mux_module mux_module_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3975]),.i2(intermediate_reg_0[3974]),.o(intermediate_reg_1[1987]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3973]),.i2(intermediate_reg_0[3972]),.o(intermediate_reg_1[1986]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3971]),.i2(intermediate_reg_0[3970]),.o(intermediate_reg_1[1985])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3969]),.i2(intermediate_reg_0[3968]),.o(intermediate_reg_1[1984])); 
mux_module mux_module_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3967]),.i2(intermediate_reg_0[3966]),.o(intermediate_reg_1[1983]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3965]),.i2(intermediate_reg_0[3964]),.o(intermediate_reg_1[1982])); 
mux_module mux_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3963]),.i2(intermediate_reg_0[3962]),.o(intermediate_reg_1[1981]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3961]),.i2(intermediate_reg_0[3960]),.o(intermediate_reg_1[1980])); 
fsm fsm_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3959]),.i2(intermediate_reg_0[3958]),.o(intermediate_reg_1[1979])); 
fsm fsm_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3957]),.i2(intermediate_reg_0[3956]),.o(intermediate_reg_1[1978])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3955]),.i2(intermediate_reg_0[3954]),.o(intermediate_reg_1[1977]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3953]),.i2(intermediate_reg_0[3952]),.o(intermediate_reg_1[1976]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3951]),.i2(intermediate_reg_0[3950]),.o(intermediate_reg_1[1975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3949]),.i2(intermediate_reg_0[3948]),.o(intermediate_reg_1[1974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3947]),.i2(intermediate_reg_0[3946]),.o(intermediate_reg_1[1973]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3945]),.i2(intermediate_reg_0[3944]),.o(intermediate_reg_1[1972])); 
mux_module mux_module_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3943]),.i2(intermediate_reg_0[3942]),.o(intermediate_reg_1[1971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3941]),.i2(intermediate_reg_0[3940]),.o(intermediate_reg_1[1970]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3939]),.i2(intermediate_reg_0[3938]),.o(intermediate_reg_1[1969])); 
fsm fsm_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3937]),.i2(intermediate_reg_0[3936]),.o(intermediate_reg_1[1968])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3935]),.i2(intermediate_reg_0[3934]),.o(intermediate_reg_1[1967]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3933]),.i2(intermediate_reg_0[3932]),.o(intermediate_reg_1[1966])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3931]),.i2(intermediate_reg_0[3930]),.o(intermediate_reg_1[1965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3929]),.i2(intermediate_reg_0[3928]),.o(intermediate_reg_1[1964]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3927]),.i2(intermediate_reg_0[3926]),.o(intermediate_reg_1[1963]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3925]),.i2(intermediate_reg_0[3924]),.o(intermediate_reg_1[1962])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3923]),.i2(intermediate_reg_0[3922]),.o(intermediate_reg_1[1961]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3921]),.i2(intermediate_reg_0[3920]),.o(intermediate_reg_1[1960]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3919]),.i2(intermediate_reg_0[3918]),.o(intermediate_reg_1[1959])); 
fsm fsm_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3917]),.i2(intermediate_reg_0[3916]),.o(intermediate_reg_1[1958])); 
fsm fsm_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3915]),.i2(intermediate_reg_0[3914]),.o(intermediate_reg_1[1957])); 
fsm fsm_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3913]),.i2(intermediate_reg_0[3912]),.o(intermediate_reg_1[1956])); 
mux_module mux_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3911]),.i2(intermediate_reg_0[3910]),.o(intermediate_reg_1[1955]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3909]),.i2(intermediate_reg_0[3908]),.o(intermediate_reg_1[1954]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3907]),.i2(intermediate_reg_0[3906]),.o(intermediate_reg_1[1953]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3905]),.i2(intermediate_reg_0[3904]),.o(intermediate_reg_1[1952])); 
fsm fsm_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3903]),.i2(intermediate_reg_0[3902]),.o(intermediate_reg_1[1951])); 
mux_module mux_module_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3901]),.i2(intermediate_reg_0[3900]),.o(intermediate_reg_1[1950]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3899]),.i2(intermediate_reg_0[3898]),.o(intermediate_reg_1[1949])); 
mux_module mux_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3897]),.i2(intermediate_reg_0[3896]),.o(intermediate_reg_1[1948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3895]),.i2(intermediate_reg_0[3894]),.o(intermediate_reg_1[1947]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3893]),.i2(intermediate_reg_0[3892]),.o(intermediate_reg_1[1946])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3891]),.i2(intermediate_reg_0[3890]),.o(intermediate_reg_1[1945])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3889]),.i2(intermediate_reg_0[3888]),.o(intermediate_reg_1[1944]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3887]),.i2(intermediate_reg_0[3886]),.o(intermediate_reg_1[1943])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3885]),.i2(intermediate_reg_0[3884]),.o(intermediate_reg_1[1942]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3883]),.i2(intermediate_reg_0[3882]),.o(intermediate_reg_1[1941])); 
fsm fsm_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3881]),.i2(intermediate_reg_0[3880]),.o(intermediate_reg_1[1940])); 
mux_module mux_module_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3879]),.i2(intermediate_reg_0[3878]),.o(intermediate_reg_1[1939]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3877]),.i2(intermediate_reg_0[3876]),.o(intermediate_reg_1[1938])); 
fsm fsm_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3875]),.i2(intermediate_reg_0[3874]),.o(intermediate_reg_1[1937])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3873]),.i2(intermediate_reg_0[3872]),.o(intermediate_reg_1[1936]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3871]),.i2(intermediate_reg_0[3870]),.o(intermediate_reg_1[1935]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3869]),.i2(intermediate_reg_0[3868]),.o(intermediate_reg_1[1934])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3867]),.i2(intermediate_reg_0[3866]),.o(intermediate_reg_1[1933])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3865]),.i2(intermediate_reg_0[3864]),.o(intermediate_reg_1[1932]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3863]),.i2(intermediate_reg_0[3862]),.o(intermediate_reg_1[1931]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3861]),.i2(intermediate_reg_0[3860]),.o(intermediate_reg_1[1930]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3859]),.i2(intermediate_reg_0[3858]),.o(intermediate_reg_1[1929])); 
mux_module mux_module_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3857]),.i2(intermediate_reg_0[3856]),.o(intermediate_reg_1[1928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3855]),.i2(intermediate_reg_0[3854]),.o(intermediate_reg_1[1927]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3853]),.i2(intermediate_reg_0[3852]),.o(intermediate_reg_1[1926]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3851]),.i2(intermediate_reg_0[3850]),.o(intermediate_reg_1[1925])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3849]),.i2(intermediate_reg_0[3848]),.o(intermediate_reg_1[1924]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3847]),.i2(intermediate_reg_0[3846]),.o(intermediate_reg_1[1923]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3845]),.i2(intermediate_reg_0[3844]),.o(intermediate_reg_1[1922])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3843]),.i2(intermediate_reg_0[3842]),.o(intermediate_reg_1[1921]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3841]),.i2(intermediate_reg_0[3840]),.o(intermediate_reg_1[1920])); 
fsm fsm_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3839]),.i2(intermediate_reg_0[3838]),.o(intermediate_reg_1[1919])); 
mux_module mux_module_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3837]),.i2(intermediate_reg_0[3836]),.o(intermediate_reg_1[1918]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3835]),.i2(intermediate_reg_0[3834]),.o(intermediate_reg_1[1917]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3833]),.i2(intermediate_reg_0[3832]),.o(intermediate_reg_1[1916])); 
mux_module mux_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3831]),.i2(intermediate_reg_0[3830]),.o(intermediate_reg_1[1915]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3829]),.i2(intermediate_reg_0[3828]),.o(intermediate_reg_1[1914]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3827]),.i2(intermediate_reg_0[3826]),.o(intermediate_reg_1[1913])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3825]),.i2(intermediate_reg_0[3824]),.o(intermediate_reg_1[1912]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3823]),.i2(intermediate_reg_0[3822]),.o(intermediate_reg_1[1911]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3821]),.i2(intermediate_reg_0[3820]),.o(intermediate_reg_1[1910])); 
fsm fsm_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3819]),.i2(intermediate_reg_0[3818]),.o(intermediate_reg_1[1909])); 
fsm fsm_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3817]),.i2(intermediate_reg_0[3816]),.o(intermediate_reg_1[1908])); 
mux_module mux_module_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3815]),.i2(intermediate_reg_0[3814]),.o(intermediate_reg_1[1907]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3813]),.i2(intermediate_reg_0[3812]),.o(intermediate_reg_1[1906]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3811]),.i2(intermediate_reg_0[3810]),.o(intermediate_reg_1[1905])); 
mux_module mux_module_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3809]),.i2(intermediate_reg_0[3808]),.o(intermediate_reg_1[1904]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3807]),.i2(intermediate_reg_0[3806]),.o(intermediate_reg_1[1903]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3805]),.i2(intermediate_reg_0[3804]),.o(intermediate_reg_1[1902]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3803]),.i2(intermediate_reg_0[3802]),.o(intermediate_reg_1[1901]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3801]),.i2(intermediate_reg_0[3800]),.o(intermediate_reg_1[1900])); 
mux_module mux_module_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3799]),.i2(intermediate_reg_0[3798]),.o(intermediate_reg_1[1899]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3797]),.i2(intermediate_reg_0[3796]),.o(intermediate_reg_1[1898]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3795]),.i2(intermediate_reg_0[3794]),.o(intermediate_reg_1[1897])); 
mux_module mux_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3793]),.i2(intermediate_reg_0[3792]),.o(intermediate_reg_1[1896]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3791]),.i2(intermediate_reg_0[3790]),.o(intermediate_reg_1[1895])); 
mux_module mux_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3789]),.i2(intermediate_reg_0[3788]),.o(intermediate_reg_1[1894]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3787]),.i2(intermediate_reg_0[3786]),.o(intermediate_reg_1[1893]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3785]),.i2(intermediate_reg_0[3784]),.o(intermediate_reg_1[1892]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3783]),.i2(intermediate_reg_0[3782]),.o(intermediate_reg_1[1891]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3781]),.i2(intermediate_reg_0[3780]),.o(intermediate_reg_1[1890])); 
fsm fsm_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3779]),.i2(intermediate_reg_0[3778]),.o(intermediate_reg_1[1889])); 
fsm fsm_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3777]),.i2(intermediate_reg_0[3776]),.o(intermediate_reg_1[1888])); 
mux_module mux_module_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3775]),.i2(intermediate_reg_0[3774]),.o(intermediate_reg_1[1887]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3773]),.i2(intermediate_reg_0[3772]),.o(intermediate_reg_1[1886]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3771]),.i2(intermediate_reg_0[3770]),.o(intermediate_reg_1[1885])); 
mux_module mux_module_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3769]),.i2(intermediate_reg_0[3768]),.o(intermediate_reg_1[1884]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3767]),.i2(intermediate_reg_0[3766]),.o(intermediate_reg_1[1883])); 
fsm fsm_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3765]),.i2(intermediate_reg_0[3764]),.o(intermediate_reg_1[1882])); 
mux_module mux_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3763]),.i2(intermediate_reg_0[3762]),.o(intermediate_reg_1[1881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3761]),.i2(intermediate_reg_0[3760]),.o(intermediate_reg_1[1880]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3759]),.i2(intermediate_reg_0[3758]),.o(intermediate_reg_1[1879]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3757]),.i2(intermediate_reg_0[3756]),.o(intermediate_reg_1[1878]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3755]),.i2(intermediate_reg_0[3754]),.o(intermediate_reg_1[1877])); 
mux_module mux_module_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3753]),.i2(intermediate_reg_0[3752]),.o(intermediate_reg_1[1876]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3751]),.i2(intermediate_reg_0[3750]),.o(intermediate_reg_1[1875])); 
mux_module mux_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3749]),.i2(intermediate_reg_0[3748]),.o(intermediate_reg_1[1874]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3747]),.i2(intermediate_reg_0[3746]),.o(intermediate_reg_1[1873])); 
fsm fsm_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3745]),.i2(intermediate_reg_0[3744]),.o(intermediate_reg_1[1872])); 
mux_module mux_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3743]),.i2(intermediate_reg_0[3742]),.o(intermediate_reg_1[1871]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3741]),.i2(intermediate_reg_0[3740]),.o(intermediate_reg_1[1870])); 
mux_module mux_module_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3739]),.i2(intermediate_reg_0[3738]),.o(intermediate_reg_1[1869]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3737]),.i2(intermediate_reg_0[3736]),.o(intermediate_reg_1[1868])); 
mux_module mux_module_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3735]),.i2(intermediate_reg_0[3734]),.o(intermediate_reg_1[1867]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3733]),.i2(intermediate_reg_0[3732]),.o(intermediate_reg_1[1866]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3731]),.i2(intermediate_reg_0[3730]),.o(intermediate_reg_1[1865])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3729]),.i2(intermediate_reg_0[3728]),.o(intermediate_reg_1[1864]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3727]),.i2(intermediate_reg_0[3726]),.o(intermediate_reg_1[1863]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3725]),.i2(intermediate_reg_0[3724]),.o(intermediate_reg_1[1862]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3723]),.i2(intermediate_reg_0[3722]),.o(intermediate_reg_1[1861])); 
mux_module mux_module_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3721]),.i2(intermediate_reg_0[3720]),.o(intermediate_reg_1[1860]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3719]),.i2(intermediate_reg_0[3718]),.o(intermediate_reg_1[1859])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3717]),.i2(intermediate_reg_0[3716]),.o(intermediate_reg_1[1858]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3715]),.i2(intermediate_reg_0[3714]),.o(intermediate_reg_1[1857]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3713]),.i2(intermediate_reg_0[3712]),.o(intermediate_reg_1[1856])); 
fsm fsm_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3711]),.i2(intermediate_reg_0[3710]),.o(intermediate_reg_1[1855])); 
mux_module mux_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3709]),.i2(intermediate_reg_0[3708]),.o(intermediate_reg_1[1854]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3707]),.i2(intermediate_reg_0[3706]),.o(intermediate_reg_1[1853])); 
mux_module mux_module_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3705]),.i2(intermediate_reg_0[3704]),.o(intermediate_reg_1[1852]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3703]),.i2(intermediate_reg_0[3702]),.o(intermediate_reg_1[1851])); 
fsm fsm_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3701]),.i2(intermediate_reg_0[3700]),.o(intermediate_reg_1[1850])); 
fsm fsm_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3699]),.i2(intermediate_reg_0[3698]),.o(intermediate_reg_1[1849])); 
mux_module mux_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3697]),.i2(intermediate_reg_0[3696]),.o(intermediate_reg_1[1848]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3695]),.i2(intermediate_reg_0[3694]),.o(intermediate_reg_1[1847])); 
fsm fsm_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3693]),.i2(intermediate_reg_0[3692]),.o(intermediate_reg_1[1846])); 
mux_module mux_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3691]),.i2(intermediate_reg_0[3690]),.o(intermediate_reg_1[1845]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3689]),.i2(intermediate_reg_0[3688]),.o(intermediate_reg_1[1844])); 
mux_module mux_module_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3687]),.i2(intermediate_reg_0[3686]),.o(intermediate_reg_1[1843]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3685]),.i2(intermediate_reg_0[3684]),.o(intermediate_reg_1[1842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3683]),.i2(intermediate_reg_0[3682]),.o(intermediate_reg_1[1841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3681]),.i2(intermediate_reg_0[3680]),.o(intermediate_reg_1[1840]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3679]),.i2(intermediate_reg_0[3678]),.o(intermediate_reg_1[1839]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3677]),.i2(intermediate_reg_0[3676]),.o(intermediate_reg_1[1838])); 
fsm fsm_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3675]),.i2(intermediate_reg_0[3674]),.o(intermediate_reg_1[1837])); 
fsm fsm_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3673]),.i2(intermediate_reg_0[3672]),.o(intermediate_reg_1[1836])); 
fsm fsm_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3671]),.i2(intermediate_reg_0[3670]),.o(intermediate_reg_1[1835])); 
fsm fsm_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3669]),.i2(intermediate_reg_0[3668]),.o(intermediate_reg_1[1834])); 
fsm fsm_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3667]),.i2(intermediate_reg_0[3666]),.o(intermediate_reg_1[1833])); 
fsm fsm_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3665]),.i2(intermediate_reg_0[3664]),.o(intermediate_reg_1[1832])); 
fsm fsm_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3663]),.i2(intermediate_reg_0[3662]),.o(intermediate_reg_1[1831])); 
fsm fsm_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3661]),.i2(intermediate_reg_0[3660]),.o(intermediate_reg_1[1830])); 
mux_module mux_module_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3659]),.i2(intermediate_reg_0[3658]),.o(intermediate_reg_1[1829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3657]),.i2(intermediate_reg_0[3656]),.o(intermediate_reg_1[1828]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3655]),.i2(intermediate_reg_0[3654]),.o(intermediate_reg_1[1827])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3653]),.i2(intermediate_reg_0[3652]),.o(intermediate_reg_1[1826])); 
fsm fsm_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3651]),.i2(intermediate_reg_0[3650]),.o(intermediate_reg_1[1825])); 
mux_module mux_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3649]),.i2(intermediate_reg_0[3648]),.o(intermediate_reg_1[1824]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3647]),.i2(intermediate_reg_0[3646]),.o(intermediate_reg_1[1823]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3645]),.i2(intermediate_reg_0[3644]),.o(intermediate_reg_1[1822])); 
fsm fsm_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3643]),.i2(intermediate_reg_0[3642]),.o(intermediate_reg_1[1821])); 
fsm fsm_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3641]),.i2(intermediate_reg_0[3640]),.o(intermediate_reg_1[1820])); 
fsm fsm_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3639]),.i2(intermediate_reg_0[3638]),.o(intermediate_reg_1[1819])); 
mux_module mux_module_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3637]),.i2(intermediate_reg_0[3636]),.o(intermediate_reg_1[1818]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3635]),.i2(intermediate_reg_0[3634]),.o(intermediate_reg_1[1817]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3633]),.i2(intermediate_reg_0[3632]),.o(intermediate_reg_1[1816])); 
mux_module mux_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3631]),.i2(intermediate_reg_0[3630]),.o(intermediate_reg_1[1815]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3629]),.i2(intermediate_reg_0[3628]),.o(intermediate_reg_1[1814])); 
mux_module mux_module_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3627]),.i2(intermediate_reg_0[3626]),.o(intermediate_reg_1[1813]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3625]),.i2(intermediate_reg_0[3624]),.o(intermediate_reg_1[1812]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3623]),.i2(intermediate_reg_0[3622]),.o(intermediate_reg_1[1811])); 
fsm fsm_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3621]),.i2(intermediate_reg_0[3620]),.o(intermediate_reg_1[1810])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3619]),.i2(intermediate_reg_0[3618]),.o(intermediate_reg_1[1809])); 
fsm fsm_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3617]),.i2(intermediate_reg_0[3616]),.o(intermediate_reg_1[1808])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3615]),.i2(intermediate_reg_0[3614]),.o(intermediate_reg_1[1807]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3613]),.i2(intermediate_reg_0[3612]),.o(intermediate_reg_1[1806]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3611]),.i2(intermediate_reg_0[3610]),.o(intermediate_reg_1[1805])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3609]),.i2(intermediate_reg_0[3608]),.o(intermediate_reg_1[1804])); 
fsm fsm_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3607]),.i2(intermediate_reg_0[3606]),.o(intermediate_reg_1[1803])); 
mux_module mux_module_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3605]),.i2(intermediate_reg_0[3604]),.o(intermediate_reg_1[1802]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3603]),.i2(intermediate_reg_0[3602]),.o(intermediate_reg_1[1801]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3601]),.i2(intermediate_reg_0[3600]),.o(intermediate_reg_1[1800])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3599]),.i2(intermediate_reg_0[3598]),.o(intermediate_reg_1[1799]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3597]),.i2(intermediate_reg_0[3596]),.o(intermediate_reg_1[1798])); 
mux_module mux_module_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3595]),.i2(intermediate_reg_0[3594]),.o(intermediate_reg_1[1797]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3593]),.i2(intermediate_reg_0[3592]),.o(intermediate_reg_1[1796]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3591]),.i2(intermediate_reg_0[3590]),.o(intermediate_reg_1[1795])); 
mux_module mux_module_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3589]),.i2(intermediate_reg_0[3588]),.o(intermediate_reg_1[1794]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3587]),.i2(intermediate_reg_0[3586]),.o(intermediate_reg_1[1793])); 
fsm fsm_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3585]),.i2(intermediate_reg_0[3584]),.o(intermediate_reg_1[1792])); 
fsm fsm_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3583]),.i2(intermediate_reg_0[3582]),.o(intermediate_reg_1[1791])); 
fsm fsm_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3581]),.i2(intermediate_reg_0[3580]),.o(intermediate_reg_1[1790])); 
mux_module mux_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3579]),.i2(intermediate_reg_0[3578]),.o(intermediate_reg_1[1789]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3577]),.i2(intermediate_reg_0[3576]),.o(intermediate_reg_1[1788])); 
fsm fsm_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3575]),.i2(intermediate_reg_0[3574]),.o(intermediate_reg_1[1787])); 
mux_module mux_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3573]),.i2(intermediate_reg_0[3572]),.o(intermediate_reg_1[1786]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3571]),.i2(intermediate_reg_0[3570]),.o(intermediate_reg_1[1785])); 
fsm fsm_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3569]),.i2(intermediate_reg_0[3568]),.o(intermediate_reg_1[1784])); 
fsm fsm_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3567]),.i2(intermediate_reg_0[3566]),.o(intermediate_reg_1[1783])); 
mux_module mux_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3565]),.i2(intermediate_reg_0[3564]),.o(intermediate_reg_1[1782]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3563]),.i2(intermediate_reg_0[3562]),.o(intermediate_reg_1[1781]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3561]),.i2(intermediate_reg_0[3560]),.o(intermediate_reg_1[1780]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3559]),.i2(intermediate_reg_0[3558]),.o(intermediate_reg_1[1779]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3557]),.i2(intermediate_reg_0[3556]),.o(intermediate_reg_1[1778])); 
fsm fsm_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3555]),.i2(intermediate_reg_0[3554]),.o(intermediate_reg_1[1777])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3553]),.i2(intermediate_reg_0[3552]),.o(intermediate_reg_1[1776]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3551]),.i2(intermediate_reg_0[3550]),.o(intermediate_reg_1[1775])); 
fsm fsm_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3549]),.i2(intermediate_reg_0[3548]),.o(intermediate_reg_1[1774])); 
mux_module mux_module_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3547]),.i2(intermediate_reg_0[3546]),.o(intermediate_reg_1[1773]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3545]),.i2(intermediate_reg_0[3544]),.o(intermediate_reg_1[1772]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3543]),.i2(intermediate_reg_0[3542]),.o(intermediate_reg_1[1771]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3541]),.i2(intermediate_reg_0[3540]),.o(intermediate_reg_1[1770])); 
fsm fsm_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3539]),.i2(intermediate_reg_0[3538]),.o(intermediate_reg_1[1769])); 
mux_module mux_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3537]),.i2(intermediate_reg_0[3536]),.o(intermediate_reg_1[1768]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3535]),.i2(intermediate_reg_0[3534]),.o(intermediate_reg_1[1767])); 
mux_module mux_module_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3533]),.i2(intermediate_reg_0[3532]),.o(intermediate_reg_1[1766]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3531]),.i2(intermediate_reg_0[3530]),.o(intermediate_reg_1[1765])); 
fsm fsm_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3529]),.i2(intermediate_reg_0[3528]),.o(intermediate_reg_1[1764])); 
fsm fsm_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3527]),.i2(intermediate_reg_0[3526]),.o(intermediate_reg_1[1763])); 
fsm fsm_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3525]),.i2(intermediate_reg_0[3524]),.o(intermediate_reg_1[1762])); 
fsm fsm_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3523]),.i2(intermediate_reg_0[3522]),.o(intermediate_reg_1[1761])); 
mux_module mux_module_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3521]),.i2(intermediate_reg_0[3520]),.o(intermediate_reg_1[1760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3519]),.i2(intermediate_reg_0[3518]),.o(intermediate_reg_1[1759]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3517]),.i2(intermediate_reg_0[3516]),.o(intermediate_reg_1[1758])); 
fsm fsm_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3515]),.i2(intermediate_reg_0[3514]),.o(intermediate_reg_1[1757])); 
fsm fsm_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3513]),.i2(intermediate_reg_0[3512]),.o(intermediate_reg_1[1756])); 
fsm fsm_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3511]),.i2(intermediate_reg_0[3510]),.o(intermediate_reg_1[1755])); 
fsm fsm_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3509]),.i2(intermediate_reg_0[3508]),.o(intermediate_reg_1[1754])); 
fsm fsm_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3507]),.i2(intermediate_reg_0[3506]),.o(intermediate_reg_1[1753])); 
fsm fsm_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3505]),.i2(intermediate_reg_0[3504]),.o(intermediate_reg_1[1752])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3503]),.i2(intermediate_reg_0[3502]),.o(intermediate_reg_1[1751]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3501]),.i2(intermediate_reg_0[3500]),.o(intermediate_reg_1[1750]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3499]),.i2(intermediate_reg_0[3498]),.o(intermediate_reg_1[1749])); 
mux_module mux_module_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3497]),.i2(intermediate_reg_0[3496]),.o(intermediate_reg_1[1748]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3495]),.i2(intermediate_reg_0[3494]),.o(intermediate_reg_1[1747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3493]),.i2(intermediate_reg_0[3492]),.o(intermediate_reg_1[1746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3491]),.i2(intermediate_reg_0[3490]),.o(intermediate_reg_1[1745]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3489]),.i2(intermediate_reg_0[3488]),.o(intermediate_reg_1[1744])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3487]),.i2(intermediate_reg_0[3486]),.o(intermediate_reg_1[1743]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3485]),.i2(intermediate_reg_0[3484]),.o(intermediate_reg_1[1742])); 
fsm fsm_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3483]),.i2(intermediate_reg_0[3482]),.o(intermediate_reg_1[1741])); 
fsm fsm_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3481]),.i2(intermediate_reg_0[3480]),.o(intermediate_reg_1[1740])); 
fsm fsm_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3479]),.i2(intermediate_reg_0[3478]),.o(intermediate_reg_1[1739])); 
mux_module mux_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3477]),.i2(intermediate_reg_0[3476]),.o(intermediate_reg_1[1738]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3475]),.i2(intermediate_reg_0[3474]),.o(intermediate_reg_1[1737])); 
mux_module mux_module_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3473]),.i2(intermediate_reg_0[3472]),.o(intermediate_reg_1[1736]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3471]),.i2(intermediate_reg_0[3470]),.o(intermediate_reg_1[1735])); 
fsm fsm_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3469]),.i2(intermediate_reg_0[3468]),.o(intermediate_reg_1[1734])); 
fsm fsm_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3467]),.i2(intermediate_reg_0[3466]),.o(intermediate_reg_1[1733])); 
fsm fsm_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3465]),.i2(intermediate_reg_0[3464]),.o(intermediate_reg_1[1732])); 
mux_module mux_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3463]),.i2(intermediate_reg_0[3462]),.o(intermediate_reg_1[1731]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3461]),.i2(intermediate_reg_0[3460]),.o(intermediate_reg_1[1730]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3459]),.i2(intermediate_reg_0[3458]),.o(intermediate_reg_1[1729]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3457]),.i2(intermediate_reg_0[3456]),.o(intermediate_reg_1[1728])); 
fsm fsm_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3455]),.i2(intermediate_reg_0[3454]),.o(intermediate_reg_1[1727])); 
fsm fsm_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3453]),.i2(intermediate_reg_0[3452]),.o(intermediate_reg_1[1726])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3451]),.i2(intermediate_reg_0[3450]),.o(intermediate_reg_1[1725])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3449]),.i2(intermediate_reg_0[3448]),.o(intermediate_reg_1[1724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3447]),.i2(intermediate_reg_0[3446]),.o(intermediate_reg_1[1723]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3445]),.i2(intermediate_reg_0[3444]),.o(intermediate_reg_1[1722]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3443]),.i2(intermediate_reg_0[3442]),.o(intermediate_reg_1[1721]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3441]),.i2(intermediate_reg_0[3440]),.o(intermediate_reg_1[1720]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3439]),.i2(intermediate_reg_0[3438]),.o(intermediate_reg_1[1719]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3437]),.i2(intermediate_reg_0[3436]),.o(intermediate_reg_1[1718])); 
mux_module mux_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3435]),.i2(intermediate_reg_0[3434]),.o(intermediate_reg_1[1717]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3433]),.i2(intermediate_reg_0[3432]),.o(intermediate_reg_1[1716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3431]),.i2(intermediate_reg_0[3430]),.o(intermediate_reg_1[1715]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3429]),.i2(intermediate_reg_0[3428]),.o(intermediate_reg_1[1714])); 
mux_module mux_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3427]),.i2(intermediate_reg_0[3426]),.o(intermediate_reg_1[1713]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3425]),.i2(intermediate_reg_0[3424]),.o(intermediate_reg_1[1712])); 
mux_module mux_module_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3423]),.i2(intermediate_reg_0[3422]),.o(intermediate_reg_1[1711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3421]),.i2(intermediate_reg_0[3420]),.o(intermediate_reg_1[1710]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3419]),.i2(intermediate_reg_0[3418]),.o(intermediate_reg_1[1709]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3417]),.i2(intermediate_reg_0[3416]),.o(intermediate_reg_1[1708]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3415]),.i2(intermediate_reg_0[3414]),.o(intermediate_reg_1[1707])); 
fsm fsm_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3413]),.i2(intermediate_reg_0[3412]),.o(intermediate_reg_1[1706])); 
fsm fsm_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3411]),.i2(intermediate_reg_0[3410]),.o(intermediate_reg_1[1705])); 
fsm fsm_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3409]),.i2(intermediate_reg_0[3408]),.o(intermediate_reg_1[1704])); 
mux_module mux_module_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3407]),.i2(intermediate_reg_0[3406]),.o(intermediate_reg_1[1703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3405]),.i2(intermediate_reg_0[3404]),.o(intermediate_reg_1[1702]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3403]),.i2(intermediate_reg_0[3402]),.o(intermediate_reg_1[1701])); 
mux_module mux_module_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3401]),.i2(intermediate_reg_0[3400]),.o(intermediate_reg_1[1700]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3399]),.i2(intermediate_reg_0[3398]),.o(intermediate_reg_1[1699]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3397]),.i2(intermediate_reg_0[3396]),.o(intermediate_reg_1[1698])); 
fsm fsm_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3395]),.i2(intermediate_reg_0[3394]),.o(intermediate_reg_1[1697])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3393]),.i2(intermediate_reg_0[3392]),.o(intermediate_reg_1[1696]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3391]),.i2(intermediate_reg_0[3390]),.o(intermediate_reg_1[1695])); 
mux_module mux_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3389]),.i2(intermediate_reg_0[3388]),.o(intermediate_reg_1[1694]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3387]),.i2(intermediate_reg_0[3386]),.o(intermediate_reg_1[1693])); 
mux_module mux_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3385]),.i2(intermediate_reg_0[3384]),.o(intermediate_reg_1[1692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3383]),.i2(intermediate_reg_0[3382]),.o(intermediate_reg_1[1691]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3381]),.i2(intermediate_reg_0[3380]),.o(intermediate_reg_1[1690]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3379]),.i2(intermediate_reg_0[3378]),.o(intermediate_reg_1[1689])); 
mux_module mux_module_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3377]),.i2(intermediate_reg_0[3376]),.o(intermediate_reg_1[1688]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3375]),.i2(intermediate_reg_0[3374]),.o(intermediate_reg_1[1687])); 
fsm fsm_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3373]),.i2(intermediate_reg_0[3372]),.o(intermediate_reg_1[1686])); 
fsm fsm_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3371]),.i2(intermediate_reg_0[3370]),.o(intermediate_reg_1[1685])); 
fsm fsm_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3369]),.i2(intermediate_reg_0[3368]),.o(intermediate_reg_1[1684])); 
fsm fsm_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3367]),.i2(intermediate_reg_0[3366]),.o(intermediate_reg_1[1683])); 
fsm fsm_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3365]),.i2(intermediate_reg_0[3364]),.o(intermediate_reg_1[1682])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3363]),.i2(intermediate_reg_0[3362]),.o(intermediate_reg_1[1681])); 
mux_module mux_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3361]),.i2(intermediate_reg_0[3360]),.o(intermediate_reg_1[1680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3359]),.i2(intermediate_reg_0[3358]),.o(intermediate_reg_1[1679]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3357]),.i2(intermediate_reg_0[3356]),.o(intermediate_reg_1[1678])); 
mux_module mux_module_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3355]),.i2(intermediate_reg_0[3354]),.o(intermediate_reg_1[1677]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3353]),.i2(intermediate_reg_0[3352]),.o(intermediate_reg_1[1676])); 
mux_module mux_module_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3351]),.i2(intermediate_reg_0[3350]),.o(intermediate_reg_1[1675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3349]),.i2(intermediate_reg_0[3348]),.o(intermediate_reg_1[1674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3347]),.i2(intermediate_reg_0[3346]),.o(intermediate_reg_1[1673]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3345]),.i2(intermediate_reg_0[3344]),.o(intermediate_reg_1[1672]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3343]),.i2(intermediate_reg_0[3342]),.o(intermediate_reg_1[1671])); 
mux_module mux_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3341]),.i2(intermediate_reg_0[3340]),.o(intermediate_reg_1[1670]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3339]),.i2(intermediate_reg_0[3338]),.o(intermediate_reg_1[1669]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3337]),.i2(intermediate_reg_0[3336]),.o(intermediate_reg_1[1668])); 
fsm fsm_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3335]),.i2(intermediate_reg_0[3334]),.o(intermediate_reg_1[1667])); 
fsm fsm_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3333]),.i2(intermediate_reg_0[3332]),.o(intermediate_reg_1[1666])); 
fsm fsm_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3331]),.i2(intermediate_reg_0[3330]),.o(intermediate_reg_1[1665])); 
fsm fsm_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3329]),.i2(intermediate_reg_0[3328]),.o(intermediate_reg_1[1664])); 
mux_module mux_module_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3327]),.i2(intermediate_reg_0[3326]),.o(intermediate_reg_1[1663]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3325]),.i2(intermediate_reg_0[3324]),.o(intermediate_reg_1[1662]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3323]),.i2(intermediate_reg_0[3322]),.o(intermediate_reg_1[1661]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3321]),.i2(intermediate_reg_0[3320]),.o(intermediate_reg_1[1660]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3319]),.i2(intermediate_reg_0[3318]),.o(intermediate_reg_1[1659])); 
mux_module mux_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3317]),.i2(intermediate_reg_0[3316]),.o(intermediate_reg_1[1658]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3315]),.i2(intermediate_reg_0[3314]),.o(intermediate_reg_1[1657])); 
mux_module mux_module_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3313]),.i2(intermediate_reg_0[3312]),.o(intermediate_reg_1[1656]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3311]),.i2(intermediate_reg_0[3310]),.o(intermediate_reg_1[1655])); 
fsm fsm_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3309]),.i2(intermediate_reg_0[3308]),.o(intermediate_reg_1[1654])); 
mux_module mux_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3307]),.i2(intermediate_reg_0[3306]),.o(intermediate_reg_1[1653]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3305]),.i2(intermediate_reg_0[3304]),.o(intermediate_reg_1[1652]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3303]),.i2(intermediate_reg_0[3302]),.o(intermediate_reg_1[1651])); 
mux_module mux_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3301]),.i2(intermediate_reg_0[3300]),.o(intermediate_reg_1[1650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3299]),.i2(intermediate_reg_0[3298]),.o(intermediate_reg_1[1649]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3297]),.i2(intermediate_reg_0[3296]),.o(intermediate_reg_1[1648])); 
mux_module mux_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3295]),.i2(intermediate_reg_0[3294]),.o(intermediate_reg_1[1647]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3293]),.i2(intermediate_reg_0[3292]),.o(intermediate_reg_1[1646])); 
mux_module mux_module_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3291]),.i2(intermediate_reg_0[3290]),.o(intermediate_reg_1[1645]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3289]),.i2(intermediate_reg_0[3288]),.o(intermediate_reg_1[1644])); 
fsm fsm_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3287]),.i2(intermediate_reg_0[3286]),.o(intermediate_reg_1[1643])); 
mux_module mux_module_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3285]),.i2(intermediate_reg_0[3284]),.o(intermediate_reg_1[1642]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3283]),.i2(intermediate_reg_0[3282]),.o(intermediate_reg_1[1641]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3281]),.i2(intermediate_reg_0[3280]),.o(intermediate_reg_1[1640]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3279]),.i2(intermediate_reg_0[3278]),.o(intermediate_reg_1[1639]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3277]),.i2(intermediate_reg_0[3276]),.o(intermediate_reg_1[1638])); 
fsm fsm_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3275]),.i2(intermediate_reg_0[3274]),.o(intermediate_reg_1[1637])); 
mux_module mux_module_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3273]),.i2(intermediate_reg_0[3272]),.o(intermediate_reg_1[1636]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3271]),.i2(intermediate_reg_0[3270]),.o(intermediate_reg_1[1635]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3269]),.i2(intermediate_reg_0[3268]),.o(intermediate_reg_1[1634]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3267]),.i2(intermediate_reg_0[3266]),.o(intermediate_reg_1[1633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3265]),.i2(intermediate_reg_0[3264]),.o(intermediate_reg_1[1632]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3263]),.i2(intermediate_reg_0[3262]),.o(intermediate_reg_1[1631]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3261]),.i2(intermediate_reg_0[3260]),.o(intermediate_reg_1[1630]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3259]),.i2(intermediate_reg_0[3258]),.o(intermediate_reg_1[1629])); 
mux_module mux_module_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3257]),.i2(intermediate_reg_0[3256]),.o(intermediate_reg_1[1628]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3255]),.i2(intermediate_reg_0[3254]),.o(intermediate_reg_1[1627])); 
mux_module mux_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3253]),.i2(intermediate_reg_0[3252]),.o(intermediate_reg_1[1626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3251]),.i2(intermediate_reg_0[3250]),.o(intermediate_reg_1[1625])); 
mux_module mux_module_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3249]),.i2(intermediate_reg_0[3248]),.o(intermediate_reg_1[1624]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3247]),.i2(intermediate_reg_0[3246]),.o(intermediate_reg_1[1623])); 
fsm fsm_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3245]),.i2(intermediate_reg_0[3244]),.o(intermediate_reg_1[1622])); 
mux_module mux_module_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3243]),.i2(intermediate_reg_0[3242]),.o(intermediate_reg_1[1621]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3241]),.i2(intermediate_reg_0[3240]),.o(intermediate_reg_1[1620]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3239]),.i2(intermediate_reg_0[3238]),.o(intermediate_reg_1[1619])); 
fsm fsm_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3237]),.i2(intermediate_reg_0[3236]),.o(intermediate_reg_1[1618])); 
fsm fsm_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3235]),.i2(intermediate_reg_0[3234]),.o(intermediate_reg_1[1617])); 
fsm fsm_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3233]),.i2(intermediate_reg_0[3232]),.o(intermediate_reg_1[1616])); 
mux_module mux_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3231]),.i2(intermediate_reg_0[3230]),.o(intermediate_reg_1[1615]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3229]),.i2(intermediate_reg_0[3228]),.o(intermediate_reg_1[1614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3227]),.i2(intermediate_reg_0[3226]),.o(intermediate_reg_1[1613]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3225]),.i2(intermediate_reg_0[3224]),.o(intermediate_reg_1[1612])); 
fsm fsm_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3223]),.i2(intermediate_reg_0[3222]),.o(intermediate_reg_1[1611])); 
mux_module mux_module_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3221]),.i2(intermediate_reg_0[3220]),.o(intermediate_reg_1[1610]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3219]),.i2(intermediate_reg_0[3218]),.o(intermediate_reg_1[1609]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3217]),.i2(intermediate_reg_0[3216]),.o(intermediate_reg_1[1608])); 
mux_module mux_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3215]),.i2(intermediate_reg_0[3214]),.o(intermediate_reg_1[1607]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3213]),.i2(intermediate_reg_0[3212]),.o(intermediate_reg_1[1606])); 
mux_module mux_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3211]),.i2(intermediate_reg_0[3210]),.o(intermediate_reg_1[1605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3209]),.i2(intermediate_reg_0[3208]),.o(intermediate_reg_1[1604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3207]),.i2(intermediate_reg_0[3206]),.o(intermediate_reg_1[1603]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3205]),.i2(intermediate_reg_0[3204]),.o(intermediate_reg_1[1602])); 
fsm fsm_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3203]),.i2(intermediate_reg_0[3202]),.o(intermediate_reg_1[1601])); 
fsm fsm_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3201]),.i2(intermediate_reg_0[3200]),.o(intermediate_reg_1[1600])); 
mux_module mux_module_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3199]),.i2(intermediate_reg_0[3198]),.o(intermediate_reg_1[1599]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3197]),.i2(intermediate_reg_0[3196]),.o(intermediate_reg_1[1598])); 
mux_module mux_module_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3195]),.i2(intermediate_reg_0[3194]),.o(intermediate_reg_1[1597]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3193]),.i2(intermediate_reg_0[3192]),.o(intermediate_reg_1[1596])); 
fsm fsm_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3191]),.i2(intermediate_reg_0[3190]),.o(intermediate_reg_1[1595])); 
fsm fsm_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3189]),.i2(intermediate_reg_0[3188]),.o(intermediate_reg_1[1594])); 
fsm fsm_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3187]),.i2(intermediate_reg_0[3186]),.o(intermediate_reg_1[1593])); 
fsm fsm_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3185]),.i2(intermediate_reg_0[3184]),.o(intermediate_reg_1[1592])); 
fsm fsm_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3183]),.i2(intermediate_reg_0[3182]),.o(intermediate_reg_1[1591])); 
mux_module mux_module_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3181]),.i2(intermediate_reg_0[3180]),.o(intermediate_reg_1[1590]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3179]),.i2(intermediate_reg_0[3178]),.o(intermediate_reg_1[1589])); 
fsm fsm_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3177]),.i2(intermediate_reg_0[3176]),.o(intermediate_reg_1[1588])); 
fsm fsm_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3175]),.i2(intermediate_reg_0[3174]),.o(intermediate_reg_1[1587])); 
mux_module mux_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3173]),.i2(intermediate_reg_0[3172]),.o(intermediate_reg_1[1586]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3171]),.i2(intermediate_reg_0[3170]),.o(intermediate_reg_1[1585])); 
mux_module mux_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3169]),.i2(intermediate_reg_0[3168]),.o(intermediate_reg_1[1584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3167]),.i2(intermediate_reg_0[3166]),.o(intermediate_reg_1[1583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3165]),.i2(intermediate_reg_0[3164]),.o(intermediate_reg_1[1582]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3163]),.i2(intermediate_reg_0[3162]),.o(intermediate_reg_1[1581])); 
mux_module mux_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3161]),.i2(intermediate_reg_0[3160]),.o(intermediate_reg_1[1580]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3159]),.i2(intermediate_reg_0[3158]),.o(intermediate_reg_1[1579])); 
fsm fsm_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3157]),.i2(intermediate_reg_0[3156]),.o(intermediate_reg_1[1578])); 
fsm fsm_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3155]),.i2(intermediate_reg_0[3154]),.o(intermediate_reg_1[1577])); 
mux_module mux_module_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3153]),.i2(intermediate_reg_0[3152]),.o(intermediate_reg_1[1576]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3151]),.i2(intermediate_reg_0[3150]),.o(intermediate_reg_1[1575]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3149]),.i2(intermediate_reg_0[3148]),.o(intermediate_reg_1[1574]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3147]),.i2(intermediate_reg_0[3146]),.o(intermediate_reg_1[1573]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3145]),.i2(intermediate_reg_0[3144]),.o(intermediate_reg_1[1572])); 
mux_module mux_module_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3143]),.i2(intermediate_reg_0[3142]),.o(intermediate_reg_1[1571]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3141]),.i2(intermediate_reg_0[3140]),.o(intermediate_reg_1[1570]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3139]),.i2(intermediate_reg_0[3138]),.o(intermediate_reg_1[1569])); 
fsm fsm_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3137]),.i2(intermediate_reg_0[3136]),.o(intermediate_reg_1[1568])); 
fsm fsm_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3135]),.i2(intermediate_reg_0[3134]),.o(intermediate_reg_1[1567])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3133]),.i2(intermediate_reg_0[3132]),.o(intermediate_reg_1[1566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3131]),.i2(intermediate_reg_0[3130]),.o(intermediate_reg_1[1565]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3129]),.i2(intermediate_reg_0[3128]),.o(intermediate_reg_1[1564])); 
mux_module mux_module_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3127]),.i2(intermediate_reg_0[3126]),.o(intermediate_reg_1[1563]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3125]),.i2(intermediate_reg_0[3124]),.o(intermediate_reg_1[1562]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3123]),.i2(intermediate_reg_0[3122]),.o(intermediate_reg_1[1561])); 
mux_module mux_module_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3121]),.i2(intermediate_reg_0[3120]),.o(intermediate_reg_1[1560]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3119]),.i2(intermediate_reg_0[3118]),.o(intermediate_reg_1[1559])); 
fsm fsm_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3117]),.i2(intermediate_reg_0[3116]),.o(intermediate_reg_1[1558])); 
fsm fsm_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3115]),.i2(intermediate_reg_0[3114]),.o(intermediate_reg_1[1557])); 
mux_module mux_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3113]),.i2(intermediate_reg_0[3112]),.o(intermediate_reg_1[1556]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3111]),.i2(intermediate_reg_0[3110]),.o(intermediate_reg_1[1555])); 
mux_module mux_module_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3109]),.i2(intermediate_reg_0[3108]),.o(intermediate_reg_1[1554]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3107]),.i2(intermediate_reg_0[3106]),.o(intermediate_reg_1[1553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3105]),.i2(intermediate_reg_0[3104]),.o(intermediate_reg_1[1552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3103]),.i2(intermediate_reg_0[3102]),.o(intermediate_reg_1[1551]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3101]),.i2(intermediate_reg_0[3100]),.o(intermediate_reg_1[1550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3099]),.i2(intermediate_reg_0[3098]),.o(intermediate_reg_1[1549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3097]),.i2(intermediate_reg_0[3096]),.o(intermediate_reg_1[1548]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3095]),.i2(intermediate_reg_0[3094]),.o(intermediate_reg_1[1547])); 
fsm fsm_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3093]),.i2(intermediate_reg_0[3092]),.o(intermediate_reg_1[1546])); 
fsm fsm_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3091]),.i2(intermediate_reg_0[3090]),.o(intermediate_reg_1[1545])); 
mux_module mux_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3089]),.i2(intermediate_reg_0[3088]),.o(intermediate_reg_1[1544]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3087]),.i2(intermediate_reg_0[3086]),.o(intermediate_reg_1[1543]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3085]),.i2(intermediate_reg_0[3084]),.o(intermediate_reg_1[1542])); 
fsm fsm_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3083]),.i2(intermediate_reg_0[3082]),.o(intermediate_reg_1[1541])); 
fsm fsm_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3081]),.i2(intermediate_reg_0[3080]),.o(intermediate_reg_1[1540])); 
fsm fsm_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3079]),.i2(intermediate_reg_0[3078]),.o(intermediate_reg_1[1539])); 
fsm fsm_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3077]),.i2(intermediate_reg_0[3076]),.o(intermediate_reg_1[1538])); 
fsm fsm_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3075]),.i2(intermediate_reg_0[3074]),.o(intermediate_reg_1[1537])); 
mux_module mux_module_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3073]),.i2(intermediate_reg_0[3072]),.o(intermediate_reg_1[1536]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3071]),.i2(intermediate_reg_0[3070]),.o(intermediate_reg_1[1535]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3069]),.i2(intermediate_reg_0[3068]),.o(intermediate_reg_1[1534])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3067]),.i2(intermediate_reg_0[3066]),.o(intermediate_reg_1[1533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3065]),.i2(intermediate_reg_0[3064]),.o(intermediate_reg_1[1532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3063]),.i2(intermediate_reg_0[3062]),.o(intermediate_reg_1[1531]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3061]),.i2(intermediate_reg_0[3060]),.o(intermediate_reg_1[1530])); 
fsm fsm_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3059]),.i2(intermediate_reg_0[3058]),.o(intermediate_reg_1[1529])); 
mux_module mux_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3057]),.i2(intermediate_reg_0[3056]),.o(intermediate_reg_1[1528]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3055]),.i2(intermediate_reg_0[3054]),.o(intermediate_reg_1[1527])); 
mux_module mux_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3053]),.i2(intermediate_reg_0[3052]),.o(intermediate_reg_1[1526]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3051]),.i2(intermediate_reg_0[3050]),.o(intermediate_reg_1[1525]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3049]),.i2(intermediate_reg_0[3048]),.o(intermediate_reg_1[1524])); 
mux_module mux_module_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3047]),.i2(intermediate_reg_0[3046]),.o(intermediate_reg_1[1523]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3045]),.i2(intermediate_reg_0[3044]),.o(intermediate_reg_1[1522])); 
mux_module mux_module_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3043]),.i2(intermediate_reg_0[3042]),.o(intermediate_reg_1[1521]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3041]),.i2(intermediate_reg_0[3040]),.o(intermediate_reg_1[1520]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3039]),.i2(intermediate_reg_0[3038]),.o(intermediate_reg_1[1519])); 
fsm fsm_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3037]),.i2(intermediate_reg_0[3036]),.o(intermediate_reg_1[1518])); 
fsm fsm_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3035]),.i2(intermediate_reg_0[3034]),.o(intermediate_reg_1[1517])); 
fsm fsm_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3033]),.i2(intermediate_reg_0[3032]),.o(intermediate_reg_1[1516])); 
fsm fsm_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3031]),.i2(intermediate_reg_0[3030]),.o(intermediate_reg_1[1515])); 
fsm fsm_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3029]),.i2(intermediate_reg_0[3028]),.o(intermediate_reg_1[1514])); 
fsm fsm_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3027]),.i2(intermediate_reg_0[3026]),.o(intermediate_reg_1[1513])); 
mux_module mux_module_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3025]),.i2(intermediate_reg_0[3024]),.o(intermediate_reg_1[1512]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3023]),.i2(intermediate_reg_0[3022]),.o(intermediate_reg_1[1511])); 
fsm fsm_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3021]),.i2(intermediate_reg_0[3020]),.o(intermediate_reg_1[1510])); 
mux_module mux_module_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3019]),.i2(intermediate_reg_0[3018]),.o(intermediate_reg_1[1509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3017]),.i2(intermediate_reg_0[3016]),.o(intermediate_reg_1[1508]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3015]),.i2(intermediate_reg_0[3014]),.o(intermediate_reg_1[1507]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3013]),.i2(intermediate_reg_0[3012]),.o(intermediate_reg_1[1506]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3011]),.i2(intermediate_reg_0[3010]),.o(intermediate_reg_1[1505])); 
fsm fsm_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3009]),.i2(intermediate_reg_0[3008]),.o(intermediate_reg_1[1504])); 
fsm fsm_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3007]),.i2(intermediate_reg_0[3006]),.o(intermediate_reg_1[1503])); 
mux_module mux_module_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3005]),.i2(intermediate_reg_0[3004]),.o(intermediate_reg_1[1502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3003]),.i2(intermediate_reg_0[3002]),.o(intermediate_reg_1[1501]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3001]),.i2(intermediate_reg_0[3000]),.o(intermediate_reg_1[1500])); 
fsm fsm_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2999]),.i2(intermediate_reg_0[2998]),.o(intermediate_reg_1[1499])); 
mux_module mux_module_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2997]),.i2(intermediate_reg_0[2996]),.o(intermediate_reg_1[1498]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2995]),.i2(intermediate_reg_0[2994]),.o(intermediate_reg_1[1497])); 
fsm fsm_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2993]),.i2(intermediate_reg_0[2992]),.o(intermediate_reg_1[1496])); 
fsm fsm_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2991]),.i2(intermediate_reg_0[2990]),.o(intermediate_reg_1[1495])); 
fsm fsm_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2989]),.i2(intermediate_reg_0[2988]),.o(intermediate_reg_1[1494])); 
fsm fsm_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2987]),.i2(intermediate_reg_0[2986]),.o(intermediate_reg_1[1493])); 
mux_module mux_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2985]),.i2(intermediate_reg_0[2984]),.o(intermediate_reg_1[1492]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2983]),.i2(intermediate_reg_0[2982]),.o(intermediate_reg_1[1491]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2981]),.i2(intermediate_reg_0[2980]),.o(intermediate_reg_1[1490])); 
fsm fsm_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2979]),.i2(intermediate_reg_0[2978]),.o(intermediate_reg_1[1489])); 
fsm fsm_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2977]),.i2(intermediate_reg_0[2976]),.o(intermediate_reg_1[1488])); 
fsm fsm_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2975]),.i2(intermediate_reg_0[2974]),.o(intermediate_reg_1[1487])); 
fsm fsm_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2973]),.i2(intermediate_reg_0[2972]),.o(intermediate_reg_1[1486])); 
mux_module mux_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2971]),.i2(intermediate_reg_0[2970]),.o(intermediate_reg_1[1485]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2969]),.i2(intermediate_reg_0[2968]),.o(intermediate_reg_1[1484]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2967]),.i2(intermediate_reg_0[2966]),.o(intermediate_reg_1[1483])); 
mux_module mux_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2965]),.i2(intermediate_reg_0[2964]),.o(intermediate_reg_1[1482]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2963]),.i2(intermediate_reg_0[2962]),.o(intermediate_reg_1[1481]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2961]),.i2(intermediate_reg_0[2960]),.o(intermediate_reg_1[1480])); 
mux_module mux_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2959]),.i2(intermediate_reg_0[2958]),.o(intermediate_reg_1[1479]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2957]),.i2(intermediate_reg_0[2956]),.o(intermediate_reg_1[1478])); 
mux_module mux_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2955]),.i2(intermediate_reg_0[2954]),.o(intermediate_reg_1[1477]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2953]),.i2(intermediate_reg_0[2952]),.o(intermediate_reg_1[1476])); 
fsm fsm_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2951]),.i2(intermediate_reg_0[2950]),.o(intermediate_reg_1[1475])); 
fsm fsm_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2949]),.i2(intermediate_reg_0[2948]),.o(intermediate_reg_1[1474])); 
mux_module mux_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2947]),.i2(intermediate_reg_0[2946]),.o(intermediate_reg_1[1473]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2945]),.i2(intermediate_reg_0[2944]),.o(intermediate_reg_1[1472])); 
fsm fsm_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2943]),.i2(intermediate_reg_0[2942]),.o(intermediate_reg_1[1471])); 
fsm fsm_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2941]),.i2(intermediate_reg_0[2940]),.o(intermediate_reg_1[1470])); 
mux_module mux_module_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2939]),.i2(intermediate_reg_0[2938]),.o(intermediate_reg_1[1469]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2937]),.i2(intermediate_reg_0[2936]),.o(intermediate_reg_1[1468])); 
fsm fsm_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2935]),.i2(intermediate_reg_0[2934]),.o(intermediate_reg_1[1467])); 
fsm fsm_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2933]),.i2(intermediate_reg_0[2932]),.o(intermediate_reg_1[1466])); 
fsm fsm_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2931]),.i2(intermediate_reg_0[2930]),.o(intermediate_reg_1[1465])); 
fsm fsm_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2929]),.i2(intermediate_reg_0[2928]),.o(intermediate_reg_1[1464])); 
fsm fsm_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2927]),.i2(intermediate_reg_0[2926]),.o(intermediate_reg_1[1463])); 
mux_module mux_module_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2925]),.i2(intermediate_reg_0[2924]),.o(intermediate_reg_1[1462]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2923]),.i2(intermediate_reg_0[2922]),.o(intermediate_reg_1[1461])); 
mux_module mux_module_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2921]),.i2(intermediate_reg_0[2920]),.o(intermediate_reg_1[1460]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2919]),.i2(intermediate_reg_0[2918]),.o(intermediate_reg_1[1459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2917]),.i2(intermediate_reg_0[2916]),.o(intermediate_reg_1[1458]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2915]),.i2(intermediate_reg_0[2914]),.o(intermediate_reg_1[1457]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2913]),.i2(intermediate_reg_0[2912]),.o(intermediate_reg_1[1456]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2911]),.i2(intermediate_reg_0[2910]),.o(intermediate_reg_1[1455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2909]),.i2(intermediate_reg_0[2908]),.o(intermediate_reg_1[1454]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2907]),.i2(intermediate_reg_0[2906]),.o(intermediate_reg_1[1453])); 
mux_module mux_module_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2905]),.i2(intermediate_reg_0[2904]),.o(intermediate_reg_1[1452]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2903]),.i2(intermediate_reg_0[2902]),.o(intermediate_reg_1[1451])); 
fsm fsm_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2901]),.i2(intermediate_reg_0[2900]),.o(intermediate_reg_1[1450])); 
mux_module mux_module_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2899]),.i2(intermediate_reg_0[2898]),.o(intermediate_reg_1[1449]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2897]),.i2(intermediate_reg_0[2896]),.o(intermediate_reg_1[1448])); 
fsm fsm_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2895]),.i2(intermediate_reg_0[2894]),.o(intermediate_reg_1[1447])); 
fsm fsm_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2893]),.i2(intermediate_reg_0[2892]),.o(intermediate_reg_1[1446])); 
fsm fsm_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2891]),.i2(intermediate_reg_0[2890]),.o(intermediate_reg_1[1445])); 
mux_module mux_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2889]),.i2(intermediate_reg_0[2888]),.o(intermediate_reg_1[1444]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2887]),.i2(intermediate_reg_0[2886]),.o(intermediate_reg_1[1443])); 
fsm fsm_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2885]),.i2(intermediate_reg_0[2884]),.o(intermediate_reg_1[1442])); 
mux_module mux_module_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2883]),.i2(intermediate_reg_0[2882]),.o(intermediate_reg_1[1441]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2881]),.i2(intermediate_reg_0[2880]),.o(intermediate_reg_1[1440]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2879]),.i2(intermediate_reg_0[2878]),.o(intermediate_reg_1[1439])); 
mux_module mux_module_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2877]),.i2(intermediate_reg_0[2876]),.o(intermediate_reg_1[1438]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2875]),.i2(intermediate_reg_0[2874]),.o(intermediate_reg_1[1437])); 
mux_module mux_module_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2873]),.i2(intermediate_reg_0[2872]),.o(intermediate_reg_1[1436]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2871]),.i2(intermediate_reg_0[2870]),.o(intermediate_reg_1[1435]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2869]),.i2(intermediate_reg_0[2868]),.o(intermediate_reg_1[1434])); 
mux_module mux_module_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2867]),.i2(intermediate_reg_0[2866]),.o(intermediate_reg_1[1433]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2865]),.i2(intermediate_reg_0[2864]),.o(intermediate_reg_1[1432]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2863]),.i2(intermediate_reg_0[2862]),.o(intermediate_reg_1[1431]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2861]),.i2(intermediate_reg_0[2860]),.o(intermediate_reg_1[1430])); 
fsm fsm_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2859]),.i2(intermediate_reg_0[2858]),.o(intermediate_reg_1[1429])); 
mux_module mux_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2857]),.i2(intermediate_reg_0[2856]),.o(intermediate_reg_1[1428]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2855]),.i2(intermediate_reg_0[2854]),.o(intermediate_reg_1[1427]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2853]),.i2(intermediate_reg_0[2852]),.o(intermediate_reg_1[1426])); 
mux_module mux_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2851]),.i2(intermediate_reg_0[2850]),.o(intermediate_reg_1[1425]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2849]),.i2(intermediate_reg_0[2848]),.o(intermediate_reg_1[1424]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2847]),.i2(intermediate_reg_0[2846]),.o(intermediate_reg_1[1423])); 
fsm fsm_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2845]),.i2(intermediate_reg_0[2844]),.o(intermediate_reg_1[1422])); 
fsm fsm_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2843]),.i2(intermediate_reg_0[2842]),.o(intermediate_reg_1[1421])); 
mux_module mux_module_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2841]),.i2(intermediate_reg_0[2840]),.o(intermediate_reg_1[1420]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2839]),.i2(intermediate_reg_0[2838]),.o(intermediate_reg_1[1419]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2837]),.i2(intermediate_reg_0[2836]),.o(intermediate_reg_1[1418])); 
fsm fsm_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2835]),.i2(intermediate_reg_0[2834]),.o(intermediate_reg_1[1417])); 
mux_module mux_module_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2833]),.i2(intermediate_reg_0[2832]),.o(intermediate_reg_1[1416]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2831]),.i2(intermediate_reg_0[2830]),.o(intermediate_reg_1[1415]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2829]),.i2(intermediate_reg_0[2828]),.o(intermediate_reg_1[1414]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2827]),.i2(intermediate_reg_0[2826]),.o(intermediate_reg_1[1413])); 
mux_module mux_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2825]),.i2(intermediate_reg_0[2824]),.o(intermediate_reg_1[1412]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2823]),.i2(intermediate_reg_0[2822]),.o(intermediate_reg_1[1411])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2821]),.i2(intermediate_reg_0[2820]),.o(intermediate_reg_1[1410]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2819]),.i2(intermediate_reg_0[2818]),.o(intermediate_reg_1[1409])); 
fsm fsm_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2817]),.i2(intermediate_reg_0[2816]),.o(intermediate_reg_1[1408])); 
mux_module mux_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2815]),.i2(intermediate_reg_0[2814]),.o(intermediate_reg_1[1407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2813]),.i2(intermediate_reg_0[2812]),.o(intermediate_reg_1[1406])); 
fsm fsm_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2811]),.i2(intermediate_reg_0[2810]),.o(intermediate_reg_1[1405])); 
mux_module mux_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2809]),.i2(intermediate_reg_0[2808]),.o(intermediate_reg_1[1404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2807]),.i2(intermediate_reg_0[2806]),.o(intermediate_reg_1[1403])); 
fsm fsm_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2805]),.i2(intermediate_reg_0[2804]),.o(intermediate_reg_1[1402])); 
fsm fsm_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2803]),.i2(intermediate_reg_0[2802]),.o(intermediate_reg_1[1401])); 
fsm fsm_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2801]),.i2(intermediate_reg_0[2800]),.o(intermediate_reg_1[1400])); 
fsm fsm_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2799]),.i2(intermediate_reg_0[2798]),.o(intermediate_reg_1[1399])); 
mux_module mux_module_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2797]),.i2(intermediate_reg_0[2796]),.o(intermediate_reg_1[1398]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2795]),.i2(intermediate_reg_0[2794]),.o(intermediate_reg_1[1397])); 
fsm fsm_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2793]),.i2(intermediate_reg_0[2792]),.o(intermediate_reg_1[1396])); 
fsm fsm_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2791]),.i2(intermediate_reg_0[2790]),.o(intermediate_reg_1[1395])); 
mux_module mux_module_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2789]),.i2(intermediate_reg_0[2788]),.o(intermediate_reg_1[1394]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2787]),.i2(intermediate_reg_0[2786]),.o(intermediate_reg_1[1393]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2785]),.i2(intermediate_reg_0[2784]),.o(intermediate_reg_1[1392])); 
mux_module mux_module_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2783]),.i2(intermediate_reg_0[2782]),.o(intermediate_reg_1[1391]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2781]),.i2(intermediate_reg_0[2780]),.o(intermediate_reg_1[1390])); 
mux_module mux_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2779]),.i2(intermediate_reg_0[2778]),.o(intermediate_reg_1[1389]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2777]),.i2(intermediate_reg_0[2776]),.o(intermediate_reg_1[1388]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2775]),.i2(intermediate_reg_0[2774]),.o(intermediate_reg_1[1387])); 
fsm fsm_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2773]),.i2(intermediate_reg_0[2772]),.o(intermediate_reg_1[1386])); 
mux_module mux_module_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2771]),.i2(intermediate_reg_0[2770]),.o(intermediate_reg_1[1385]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2769]),.i2(intermediate_reg_0[2768]),.o(intermediate_reg_1[1384]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2767]),.i2(intermediate_reg_0[2766]),.o(intermediate_reg_1[1383])); 
mux_module mux_module_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2765]),.i2(intermediate_reg_0[2764]),.o(intermediate_reg_1[1382]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2763]),.i2(intermediate_reg_0[2762]),.o(intermediate_reg_1[1381])); 
fsm fsm_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2761]),.i2(intermediate_reg_0[2760]),.o(intermediate_reg_1[1380])); 
fsm fsm_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2759]),.i2(intermediate_reg_0[2758]),.o(intermediate_reg_1[1379])); 
fsm fsm_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2757]),.i2(intermediate_reg_0[2756]),.o(intermediate_reg_1[1378])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2755]),.i2(intermediate_reg_0[2754]),.o(intermediate_reg_1[1377]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2753]),.i2(intermediate_reg_0[2752]),.o(intermediate_reg_1[1376])); 
fsm fsm_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2751]),.i2(intermediate_reg_0[2750]),.o(intermediate_reg_1[1375])); 
fsm fsm_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2749]),.i2(intermediate_reg_0[2748]),.o(intermediate_reg_1[1374])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2747]),.i2(intermediate_reg_0[2746]),.o(intermediate_reg_1[1373]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2745]),.i2(intermediate_reg_0[2744]),.o(intermediate_reg_1[1372])); 
mux_module mux_module_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2743]),.i2(intermediate_reg_0[2742]),.o(intermediate_reg_1[1371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2741]),.i2(intermediate_reg_0[2740]),.o(intermediate_reg_1[1370]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2739]),.i2(intermediate_reg_0[2738]),.o(intermediate_reg_1[1369]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2737]),.i2(intermediate_reg_0[2736]),.o(intermediate_reg_1[1368]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2735]),.i2(intermediate_reg_0[2734]),.o(intermediate_reg_1[1367])); 
fsm fsm_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2733]),.i2(intermediate_reg_0[2732]),.o(intermediate_reg_1[1366])); 
mux_module mux_module_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2731]),.i2(intermediate_reg_0[2730]),.o(intermediate_reg_1[1365]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2729]),.i2(intermediate_reg_0[2728]),.o(intermediate_reg_1[1364])); 
mux_module mux_module_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2727]),.i2(intermediate_reg_0[2726]),.o(intermediate_reg_1[1363]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2725]),.i2(intermediate_reg_0[2724]),.o(intermediate_reg_1[1362])); 
fsm fsm_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2723]),.i2(intermediate_reg_0[2722]),.o(intermediate_reg_1[1361])); 
mux_module mux_module_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2721]),.i2(intermediate_reg_0[2720]),.o(intermediate_reg_1[1360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2719]),.i2(intermediate_reg_0[2718]),.o(intermediate_reg_1[1359]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2717]),.i2(intermediate_reg_0[2716]),.o(intermediate_reg_1[1358])); 
fsm fsm_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2715]),.i2(intermediate_reg_0[2714]),.o(intermediate_reg_1[1357])); 
fsm fsm_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2713]),.i2(intermediate_reg_0[2712]),.o(intermediate_reg_1[1356])); 
fsm fsm_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2711]),.i2(intermediate_reg_0[2710]),.o(intermediate_reg_1[1355])); 
mux_module mux_module_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2709]),.i2(intermediate_reg_0[2708]),.o(intermediate_reg_1[1354]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2707]),.i2(intermediate_reg_0[2706]),.o(intermediate_reg_1[1353])); 
fsm fsm_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2705]),.i2(intermediate_reg_0[2704]),.o(intermediate_reg_1[1352])); 
mux_module mux_module_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2703]),.i2(intermediate_reg_0[2702]),.o(intermediate_reg_1[1351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2701]),.i2(intermediate_reg_0[2700]),.o(intermediate_reg_1[1350]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2699]),.i2(intermediate_reg_0[2698]),.o(intermediate_reg_1[1349])); 
mux_module mux_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2697]),.i2(intermediate_reg_0[2696]),.o(intermediate_reg_1[1348]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2695]),.i2(intermediate_reg_0[2694]),.o(intermediate_reg_1[1347]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2693]),.i2(intermediate_reg_0[2692]),.o(intermediate_reg_1[1346]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2691]),.i2(intermediate_reg_0[2690]),.o(intermediate_reg_1[1345])); 
mux_module mux_module_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2689]),.i2(intermediate_reg_0[2688]),.o(intermediate_reg_1[1344]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342])); 
fsm fsm_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341])); 
fsm fsm_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340])); 
fsm fsm_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339])); 
mux_module mux_module_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334])); 
fsm fsm_inst_1_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333])); 
mux_module mux_module_inst_1_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329])); 
fsm fsm_inst_1_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328])); 
fsm fsm_inst_1_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327])); 
mux_module mux_module_inst_1_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321])); 
mux_module mux_module_inst_1_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319])); 
mux_module mux_module_inst_1_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317])); 
mux_module mux_module_inst_1_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313])); 
mux_module mux_module_inst_1_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308])); 
mux_module mux_module_inst_1_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305])); 
fsm fsm_inst_1_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304])); 
fsm fsm_inst_1_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303])); 
mux_module mux_module_inst_1_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301])); 
mux_module mux_module_inst_1_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299])); 
mux_module mux_module_inst_1_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296])); 
fsm fsm_inst_1_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295])); 
mux_module mux_module_inst_1_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292])); 
fsm fsm_inst_1_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291])); 
fsm fsm_inst_1_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290])); 
fsm fsm_inst_1_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289])); 
mux_module mux_module_inst_1_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287])); 
fsm fsm_inst_1_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286])); 
fsm fsm_inst_1_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285])); 
mux_module mux_module_inst_1_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282])); 
mux_module mux_module_inst_1_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279])); 
mux_module mux_module_inst_1_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277])); 
mux_module mux_module_inst_1_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274])); 
mux_module mux_module_inst_1_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270])); 
fsm fsm_inst_1_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269])); 
fsm fsm_inst_1_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268])); 
mux_module mux_module_inst_1_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266])); 
fsm fsm_inst_1_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265])); 
fsm fsm_inst_1_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264])); 
fsm fsm_inst_1_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263])); 
mux_module mux_module_inst_1_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261])); 
mux_module mux_module_inst_1_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259])); 
mux_module mux_module_inst_1_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257])); 
fsm fsm_inst_1_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256])); 
mux_module mux_module_inst_1_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253])); 
mux_module mux_module_inst_1_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250])); 
fsm fsm_inst_1_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249])); 
mux_module mux_module_inst_1_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247])); 
fsm fsm_inst_1_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246])); 
mux_module mux_module_inst_1_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243])); 
fsm fsm_inst_1_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242])); 
mux_module mux_module_inst_1_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
mux_module mux_module_inst_1_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238])); 
fsm fsm_inst_1_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237])); 
fsm fsm_inst_1_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236])); 
fsm fsm_inst_1_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235])); 
fsm fsm_inst_1_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234])); 
mux_module mux_module_inst_1_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232])); 
mux_module mux_module_inst_1_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230])); 
mux_module mux_module_inst_1_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227])); 
mux_module mux_module_inst_1_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225])); 
mux_module mux_module_inst_1_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223])); 
fsm fsm_inst_1_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222])); 
mux_module mux_module_inst_1_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217])); 
mux_module mux_module_inst_1_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213])); 
fsm fsm_inst_1_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212])); 
fsm fsm_inst_1_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211])); 
fsm fsm_inst_1_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210])); 
mux_module mux_module_inst_1_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208])); 
fsm fsm_inst_1_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207])); 
fsm fsm_inst_1_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206])); 
mux_module mux_module_inst_1_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202])); 
mux_module mux_module_inst_1_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200])); 
mux_module mux_module_inst_1_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198])); 
mux_module mux_module_inst_1_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196])); 
fsm fsm_inst_1_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195])); 
mux_module mux_module_inst_1_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193])); 
mux_module mux_module_inst_1_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191])); 
fsm fsm_inst_1_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190])); 
fsm fsm_inst_1_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189])); 
fsm fsm_inst_1_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188])); 
mux_module mux_module_inst_1_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186])); 
fsm fsm_inst_1_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185])); 
mux_module mux_module_inst_1_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182])); 
mux_module mux_module_inst_1_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178])); 
fsm fsm_inst_1_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177])); 
fsm fsm_inst_1_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176])); 
fsm fsm_inst_1_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175])); 
mux_module mux_module_inst_1_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172])); 
fsm fsm_inst_1_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171])); 
mux_module mux_module_inst_1_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169])); 
mux_module mux_module_inst_1_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165])); 
fsm fsm_inst_1_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164])); 
mux_module mux_module_inst_1_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159])); 
mux_module mux_module_inst_1_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
fsm fsm_inst_1_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156])); 
mux_module mux_module_inst_1_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152])); 
mux_module mux_module_inst_1_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
fsm fsm_inst_1_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147])); 
mux_module mux_module_inst_1_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145])); 
mux_module mux_module_inst_1_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142])); 
mux_module mux_module_inst_1_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140])); 
fsm fsm_inst_1_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139])); 
fsm fsm_inst_1_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138])); 
fsm fsm_inst_1_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137])); 
fsm fsm_inst_1_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136])); 
fsm fsm_inst_1_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135])); 
fsm fsm_inst_1_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134])); 
mux_module mux_module_inst_1_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
mux_module mux_module_inst_1_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128])); 
fsm fsm_inst_1_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127])); 
mux_module mux_module_inst_1_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
mux_module mux_module_inst_1_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123])); 
mux_module mux_module_inst_1_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115])); 
fsm fsm_inst_1_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114])); 
mux_module mux_module_inst_1_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109])); 
fsm fsm_inst_1_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
mux_module mux_module_inst_1_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
mux_module mux_module_inst_1_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101])); 
fsm fsm_inst_1_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100])); 
mux_module mux_module_inst_1_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097])); 
fsm fsm_inst_1_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096])); 
mux_module mux_module_inst_1_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
fsm fsm_inst_1_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092])); 
fsm fsm_inst_1_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
mux_module mux_module_inst_1_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
mux_module mux_module_inst_1_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087])); 
fsm fsm_inst_1_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086])); 
fsm fsm_inst_1_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085])); 
fsm fsm_inst_1_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084])); 
fsm fsm_inst_1_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
mux_module mux_module_inst_1_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078])); 
fsm fsm_inst_1_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077])); 
fsm fsm_inst_1_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076])); 
fsm fsm_inst_1_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075])); 
fsm fsm_inst_1_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074])); 
fsm fsm_inst_1_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
fsm fsm_inst_1_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072])); 
fsm fsm_inst_1_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071])); 
mux_module mux_module_inst_1_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069])); 
mux_module mux_module_inst_1_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061])); 
fsm fsm_inst_1_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060])); 
mux_module mux_module_inst_1_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056])); 
mux_module mux_module_inst_1_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052])); 
mux_module mux_module_inst_1_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050])); 
mux_module mux_module_inst_1_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047])); 
fsm fsm_inst_1_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046])); 
mux_module mux_module_inst_1_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
fsm fsm_inst_1_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
mux_module mux_module_inst_1_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040])); 
mux_module mux_module_inst_1_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036])); 
mux_module mux_module_inst_1_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034])); 
fsm fsm_inst_1_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033])); 
mux_module mux_module_inst_1_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031])); 
mux_module mux_module_inst_1_1649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029])); 
fsm fsm_inst_1_1651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
fsm fsm_inst_1_1652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027])); 
mux_module mux_module_inst_1_1653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023])); 
mux_module mux_module_inst_1_1657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016])); 
mux_module mux_module_inst_1_1664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009])); 
mux_module mux_module_inst_1_1671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006])); 
fsm fsm_inst_1_1674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
fsm fsm_inst_1_1675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
mux_module mux_module_inst_1_1676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
mux_module mux_module_inst_1_1680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997])); 
mux_module mux_module_inst_1_1683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
mux_module mux_module_inst_1_1691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
fsm fsm_inst_1_1693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986])); 
fsm fsm_inst_1_1694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
fsm fsm_inst_1_1695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984])); 
fsm fsm_inst_1_1696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983])); 
fsm fsm_inst_1_1697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
mux_module mux_module_inst_1_1698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
fsm fsm_inst_1_1700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979])); 
mux_module mux_module_inst_1_1701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
mux_module mux_module_inst_1_1703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974])); 
mux_module mux_module_inst_1_1706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969])); 
fsm fsm_inst_1_1711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968])); 
mux_module mux_module_inst_1_1712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965])); 
fsm fsm_inst_1_1715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964])); 
mux_module mux_module_inst_1_1716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961])); 
fsm fsm_inst_1_1719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960])); 
mux_module mux_module_inst_1_1720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
mux_module mux_module_inst_1_1723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955])); 
mux_module mux_module_inst_1_1725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
fsm fsm_inst_1_1727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952])); 
fsm fsm_inst_1_1728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
mux_module mux_module_inst_1_1729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
fsm fsm_inst_1_1734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
fsm fsm_inst_1_1735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944])); 
mux_module mux_module_inst_1_1736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
mux_module mux_module_inst_1_1738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
fsm fsm_inst_1_1743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
mux_module mux_module_inst_1_1744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
mux_module mux_module_inst_1_1746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
fsm fsm_inst_1_1751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928])); 
fsm fsm_inst_1_1752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927])); 
fsm fsm_inst_1_1753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
mux_module mux_module_inst_1_1754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923])); 
mux_module mux_module_inst_1_1757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
fsm fsm_inst_1_1765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
fsm fsm_inst_1_1766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913])); 
fsm fsm_inst_1_1767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
mux_module mux_module_inst_1_1768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910])); 
fsm fsm_inst_1_1770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909])); 
mux_module mux_module_inst_1_1771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905])); 
mux_module mux_module_inst_1_1775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
fsm fsm_inst_1_1779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900])); 
fsm fsm_inst_1_1780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
mux_module mux_module_inst_1_1781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
fsm fsm_inst_1_1783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896])); 
fsm fsm_inst_1_1784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895])); 
fsm fsm_inst_1_1785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894])); 
fsm fsm_inst_1_1786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
mux_module mux_module_inst_1_1787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
mux_module mux_module_inst_1_1791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886])); 
mux_module mux_module_inst_1_1794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883])); 
fsm fsm_inst_1_1797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882])); 
mux_module mux_module_inst_1_1798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877])); 
mux_module mux_module_inst_1_1803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872])); 
fsm fsm_inst_1_1808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871])); 
fsm fsm_inst_1_1809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870])); 
mux_module mux_module_inst_1_1810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
fsm fsm_inst_1_1812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
mux_module mux_module_inst_1_1813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
mux_module mux_module_inst_1_1819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858])); 
mux_module mux_module_inst_1_1822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
fsm fsm_inst_1_1825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
mux_module mux_module_inst_1_1826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852])); 
mux_module mux_module_inst_1_1828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850])); 
fsm fsm_inst_1_1830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849])); 
mux_module mux_module_inst_1_1831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
mux_module mux_module_inst_1_1834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844])); 
fsm fsm_inst_1_1836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
mux_module mux_module_inst_1_1837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839])); 
fsm fsm_inst_1_1841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
fsm fsm_inst_1_1842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837])); 
mux_module mux_module_inst_1_1843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835])); 
fsm fsm_inst_1_1845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
fsm fsm_inst_1_1846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833])); 
mux_module mux_module_inst_1_1847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830])); 
mux_module mux_module_inst_1_1850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828])); 
fsm fsm_inst_1_1852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827])); 
fsm fsm_inst_1_1853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
mux_module mux_module_inst_1_1854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824])); 
mux_module mux_module_inst_1_1856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818])); 
mux_module mux_module_inst_1_1862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816])); 
mux_module mux_module_inst_1_1864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814])); 
fsm fsm_inst_1_1866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813])); 
fsm fsm_inst_1_1867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812])); 
fsm fsm_inst_1_1868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811])); 
mux_module mux_module_inst_1_1869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
mux_module mux_module_inst_1_1871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806])); 
fsm fsm_inst_1_1874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
fsm fsm_inst_1_1875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804])); 
mux_module mux_module_inst_1_1876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802])); 
fsm fsm_inst_1_1878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
mux_module mux_module_inst_1_1879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799])); 
fsm fsm_inst_1_1881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
mux_module mux_module_inst_1_1882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792])); 
fsm fsm_inst_1_1888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791])); 
fsm fsm_inst_1_1889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790])); 
fsm fsm_inst_1_1890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
mux_module mux_module_inst_1_1891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
fsm fsm_inst_1_1894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
mux_module mux_module_inst_1_1895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
fsm fsm_inst_1_1897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
mux_module mux_module_inst_1_1898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778])); 
mux_module mux_module_inst_1_1902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
mux_module mux_module_inst_1_1906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
mux_module mux_module_inst_1_1909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768])); 
fsm fsm_inst_1_1912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767])); 
fsm fsm_inst_1_1913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
fsm fsm_inst_1_1914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
fsm fsm_inst_1_1915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
fsm fsm_inst_1_1916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
mux_module mux_module_inst_1_1917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
fsm fsm_inst_1_1920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
mux_module mux_module_inst_1_1921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
fsm fsm_inst_1_1928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751])); 
fsm fsm_inst_1_1929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
fsm fsm_inst_1_1930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
mux_module mux_module_inst_1_1931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747])); 
fsm fsm_inst_1_1933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746])); 
fsm fsm_inst_1_1934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745])); 
fsm fsm_inst_1_1935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
fsm fsm_inst_1_1936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743])); 
mux_module mux_module_inst_1_1937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
fsm fsm_inst_1_1939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740])); 
mux_module mux_module_inst_1_1940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737])); 
fsm fsm_inst_1_1943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736])); 
mux_module mux_module_inst_1_1944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
mux_module mux_module_inst_1_1946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
mux_module mux_module_inst_1_1950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728])); 
mux_module mux_module_inst_1_1952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
mux_module mux_module_inst_1_1954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724])); 
mux_module mux_module_inst_1_1956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720])); 
mux_module mux_module_inst_1_1960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
fsm fsm_inst_1_1963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716])); 
mux_module mux_module_inst_1_1964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714])); 
fsm fsm_inst_1_1966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
fsm fsm_inst_1_1967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
mux_module mux_module_inst_1_1968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709])); 
fsm fsm_inst_1_1971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
fsm fsm_inst_1_1972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
fsm fsm_inst_1_1973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706])); 
fsm fsm_inst_1_1974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
mux_module mux_module_inst_1_1975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
mux_module mux_module_inst_1_1981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
fsm fsm_inst_1_1984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695])); 
fsm fsm_inst_1_1985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
fsm fsm_inst_1_1986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
mux_module mux_module_inst_1_1987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688])); 
mux_module mux_module_inst_1_1992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
mux_module mux_module_inst_1_1995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
fsm fsm_inst_1_1999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
fsm fsm_inst_1_2000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
fsm fsm_inst_1_2001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
mux_module mux_module_inst_1_2002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676])); 
mux_module mux_module_inst_1_2004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
mux_module mux_module_inst_1_2008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670])); 
mux_module mux_module_inst_1_2010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
mux_module mux_module_inst_1_2012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666])); 
fsm fsm_inst_1_2014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665])); 
mux_module mux_module_inst_1_2015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
mux_module mux_module_inst_1_2017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661])); 
mux_module mux_module_inst_1_2019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_2021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
fsm fsm_inst_1_2022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657])); 
fsm fsm_inst_1_2023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
fsm fsm_inst_1_2024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
mux_module mux_module_inst_1_2025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
fsm fsm_inst_1_2028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651])); 
mux_module mux_module_inst_1_2029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649])); 
fsm fsm_inst_1_2031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648])); 
fsm fsm_inst_1_2032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
mux_module mux_module_inst_1_2033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645])); 
fsm fsm_inst_1_2035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
mux_module mux_module_inst_1_2036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642])); 
fsm fsm_inst_1_2038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
mux_module mux_module_inst_1_2039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
fsm fsm_inst_1_2041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638])); 
fsm fsm_inst_1_2042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
fsm fsm_inst_1_2043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636])); 
mux_module mux_module_inst_1_2044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634])); 
mux_module mux_module_inst_1_2046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
mux_module mux_module_inst_1_2050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628])); 
fsm fsm_inst_1_2052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
mux_module mux_module_inst_1_2053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
mux_module mux_module_inst_1_2056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621])); 
mux_module mux_module_inst_1_2059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
mux_module mux_module_inst_1_2063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615])); 
fsm fsm_inst_1_2065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
mux_module mux_module_inst_1_2066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612])); 
mux_module mux_module_inst_1_2068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609])); 
fsm fsm_inst_1_2071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
mux_module mux_module_inst_1_2072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605])); 
fsm fsm_inst_1_2075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604])); 
fsm fsm_inst_1_2076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603])); 
mux_module mux_module_inst_1_2077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
fsm fsm_inst_1_2082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597])); 
mux_module mux_module_inst_1_2083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
fsm fsm_inst_1_2086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593])); 
mux_module mux_module_inst_1_2087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
mux_module mux_module_inst_1_2090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587])); 
mux_module mux_module_inst_1_2093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
fsm fsm_inst_1_2096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583])); 
mux_module mux_module_inst_1_2097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_2100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
fsm fsm_inst_1_2101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578])); 
mux_module mux_module_inst_1_2102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576])); 
mux_module mux_module_inst_1_2104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
fsm fsm_inst_1_2106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573])); 
fsm fsm_inst_1_2107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
fsm fsm_inst_1_2108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571])); 
mux_module mux_module_inst_1_2109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569])); 
mux_module mux_module_inst_1_2111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566])); 
mux_module mux_module_inst_1_2114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563])); 
fsm fsm_inst_1_2117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
fsm fsm_inst_1_2118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
mux_module mux_module_inst_1_2119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
mux_module mux_module_inst_1_2122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_2124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
mux_module mux_module_inst_1_2125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_2127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
fsm fsm_inst_1_2128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551])); 
fsm fsm_inst_1_2129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550])); 
mux_module mux_module_inst_1_2130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547])); 
mux_module mux_module_inst_1_2133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545])); 
mux_module mux_module_inst_1_2135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
fsm fsm_inst_1_2137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542])); 
fsm fsm_inst_1_2138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
mux_module mux_module_inst_1_2139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539])); 
fsm fsm_inst_1_2141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538])); 
mux_module mux_module_inst_1_2142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536])); 
fsm fsm_inst_1_2144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535])); 
fsm fsm_inst_1_2145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534])); 
mux_module mux_module_inst_1_2146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529])); 
mux_module mux_module_inst_1_2151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527])); 
mux_module mux_module_inst_1_2153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
fsm fsm_inst_1_2155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524])); 
mux_module mux_module_inst_1_2156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522])); 
fsm fsm_inst_1_2158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
fsm fsm_inst_1_2159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520])); 
mux_module mux_module_inst_1_2160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
mux_module mux_module_inst_1_2162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
fsm fsm_inst_1_2168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
mux_module mux_module_inst_1_2169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509])); 
mux_module mux_module_inst_1_2171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506])); 
fsm fsm_inst_1_2174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
fsm fsm_inst_1_2175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504])); 
mux_module mux_module_inst_1_2176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502])); 
fsm fsm_inst_1_2178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501])); 
fsm fsm_inst_1_2179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
fsm fsm_inst_1_2180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499])); 
mux_module mux_module_inst_1_2181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497])); 
mux_module mux_module_inst_1_2183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
fsm fsm_inst_1_2186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493])); 
fsm fsm_inst_1_2187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492])); 
fsm fsm_inst_1_2188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491])); 
fsm fsm_inst_1_2189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490])); 
fsm fsm_inst_1_2190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
fsm fsm_inst_1_2191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488])); 
mux_module mux_module_inst_1_2192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486])); 
fsm fsm_inst_1_2194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
mux_module mux_module_inst_1_2195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482])); 
mux_module mux_module_inst_1_2198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
fsm fsm_inst_1_2200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
fsm fsm_inst_1_2201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_2202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
mux_module mux_module_inst_1_2203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475])); 
mux_module mux_module_inst_1_2205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
fsm fsm_inst_1_2208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471])); 
fsm fsm_inst_1_2209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
mux_module mux_module_inst_1_2210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468])); 
fsm fsm_inst_1_2212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
fsm fsm_inst_1_2213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
fsm fsm_inst_1_2214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
mux_module mux_module_inst_1_2215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461])); 
fsm fsm_inst_1_2219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460])); 
fsm fsm_inst_1_2220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
fsm fsm_inst_1_2221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458])); 
mux_module mux_module_inst_1_2222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
mux_module mux_module_inst_1_2224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450])); 
fsm fsm_inst_1_2230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449])); 
fsm fsm_inst_1_2231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448])); 
mux_module mux_module_inst_1_2232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
fsm fsm_inst_1_2234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
mux_module mux_module_inst_1_2235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
fsm fsm_inst_1_2239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440])); 
fsm fsm_inst_1_2240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
fsm fsm_inst_1_2241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
fsm fsm_inst_1_2242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437])); 
mux_module mux_module_inst_1_2243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
fsm fsm_inst_1_2248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
mux_module mux_module_inst_1_2249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_2253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
mux_module mux_module_inst_1_2254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424])); 
fsm fsm_inst_1_2256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
fsm fsm_inst_1_2257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
mux_module mux_module_inst_1_2258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418])); 
mux_module mux_module_inst_1_2262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414])); 
fsm fsm_inst_1_2266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413])); 
mux_module mux_module_inst_1_2267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
fsm fsm_inst_1_2270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409])); 
mux_module mux_module_inst_1_2271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401])); 
mux_module mux_module_inst_1_2279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
mux_module mux_module_inst_1_2281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
mux_module mux_module_inst_1_2283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_2286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_2287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390])); 
fsm fsm_inst_1_2290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
mux_module mux_module_inst_1_2291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_2295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
fsm fsm_inst_1_2297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382])); 
mux_module mux_module_inst_1_2298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380])); 
mux_module mux_module_inst_1_2300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_2303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
fsm fsm_inst_1_2304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375])); 
fsm fsm_inst_1_2305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
mux_module mux_module_inst_1_2306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
fsm fsm_inst_1_2308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371])); 
mux_module mux_module_inst_1_2309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368])); 
mux_module mux_module_inst_1_2312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365])); 
mux_module mux_module_inst_1_2315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
mux_module mux_module_inst_1_2317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360])); 
mux_module mux_module_inst_1_2320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358])); 
fsm fsm_inst_1_2322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357])); 
mux_module mux_module_inst_1_2323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350])); 
mux_module mux_module_inst_1_2330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
mux_module mux_module_inst_1_2332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346])); 
fsm fsm_inst_1_2334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345])); 
fsm fsm_inst_1_2335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344])); 
mux_module mux_module_inst_1_2336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341])); 
fsm fsm_inst_1_2339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
fsm fsm_inst_1_2340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339])); 
mux_module mux_module_inst_1_2341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_2348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_2349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329])); 
fsm fsm_inst_1_2351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328])); 
fsm fsm_inst_1_2352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327])); 
mux_module mux_module_inst_1_2353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
mux_module mux_module_inst_1_2356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
mux_module mux_module_inst_1_2358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320])); 
mux_module mux_module_inst_1_2360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
mux_module mux_module_inst_1_2365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
fsm fsm_inst_1_2367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
mux_module mux_module_inst_1_2368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310])); 
mux_module mux_module_inst_1_2370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307])); 
mux_module mux_module_inst_1_2373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305])); 
mux_module mux_module_inst_1_2375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
fsm fsm_inst_1_2378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
fsm fsm_inst_1_2379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
mux_module mux_module_inst_1_2380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294])); 
mux_module mux_module_inst_1_2386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
fsm fsm_inst_1_2388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291])); 
fsm fsm_inst_1_2389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
fsm fsm_inst_1_2390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289])); 
fsm fsm_inst_1_2391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
mux_module mux_module_inst_1_2392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
mux_module mux_module_inst_1_2395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
mux_module mux_module_inst_1_2397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
fsm fsm_inst_1_2399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280])); 
mux_module mux_module_inst_1_2400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278])); 
mux_module mux_module_inst_1_2402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
fsm fsm_inst_1_2404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
mux_module mux_module_inst_1_2405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
fsm fsm_inst_1_2407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
fsm fsm_inst_1_2408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271])); 
mux_module mux_module_inst_1_2409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
fsm fsm_inst_1_2411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
fsm fsm_inst_1_2412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
mux_module mux_module_inst_1_2413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
fsm fsm_inst_1_2415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264])); 
mux_module mux_module_inst_1_2416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
fsm fsm_inst_1_2418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_2419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
fsm fsm_inst_1_2420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259])); 
fsm fsm_inst_1_2421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
fsm fsm_inst_1_2422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257])); 
mux_module mux_module_inst_1_2423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
mux_module mux_module_inst_1_2428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244])); 
mux_module mux_module_inst_1_2436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
mux_module mux_module_inst_1_2438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238])); 
mux_module mux_module_inst_1_2442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235])); 
mux_module mux_module_inst_1_2445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232])); 
mux_module mux_module_inst_1_2448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
fsm fsm_inst_1_2450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229])); 
mux_module mux_module_inst_1_2451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225])); 
mux_module mux_module_inst_1_2455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222])); 
mux_module mux_module_inst_1_2458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
mux_module mux_module_inst_1_2460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218])); 
fsm fsm_inst_1_2462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217])); 
mux_module mux_module_inst_1_2463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213])); 
mux_module mux_module_inst_1_2467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
fsm fsm_inst_1_2469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
fsm fsm_inst_1_2470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209])); 
mux_module mux_module_inst_1_2471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206])); 
fsm fsm_inst_1_2474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
fsm fsm_inst_1_2475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
mux_module mux_module_inst_1_2476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
fsm fsm_inst_1_2479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200])); 
fsm fsm_inst_1_2480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199])); 
fsm fsm_inst_1_2481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
mux_module mux_module_inst_1_2482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196])); 
mux_module mux_module_inst_1_2484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194])); 
fsm fsm_inst_1_2486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193])); 
mux_module mux_module_inst_1_2487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
mux_module mux_module_inst_1_2494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
mux_module mux_module_inst_1_2498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174])); 
fsm fsm_inst_1_2506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
mux_module mux_module_inst_1_2507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
mux_module mux_module_inst_1_2509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168])); 
mux_module mux_module_inst_1_2512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166])); 
mux_module mux_module_inst_1_2514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
mux_module mux_module_inst_1_2516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
mux_module mux_module_inst_1_2518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
fsm fsm_inst_1_2520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159])); 
mux_module mux_module_inst_1_2521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157])); 
fsm fsm_inst_1_2523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
mux_module mux_module_inst_1_2524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
mux_module mux_module_inst_1_2526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
fsm fsm_inst_1_2529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150])); 
mux_module mux_module_inst_1_2530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148])); 
mux_module mux_module_inst_1_2532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146])); 
mux_module mux_module_inst_1_2534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
mux_module mux_module_inst_1_2539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139])); 
fsm fsm_inst_1_2541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138])); 
mux_module mux_module_inst_1_2542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
fsm fsm_inst_1_2545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
fsm fsm_inst_1_2546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
fsm fsm_inst_1_2547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
fsm fsm_inst_1_2548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
fsm fsm_inst_1_2549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
fsm fsm_inst_1_2550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129])); 
fsm fsm_inst_1_2551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
fsm fsm_inst_1_2552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127])); 
fsm fsm_inst_1_2553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
fsm fsm_inst_1_2554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125])); 
fsm fsm_inst_1_2555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
mux_module mux_module_inst_1_2556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
mux_module mux_module_inst_1_2558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119])); 
fsm fsm_inst_1_2561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118])); 
mux_module mux_module_inst_1_2562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116])); 
mux_module mux_module_inst_1_2564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
fsm fsm_inst_1_2566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113])); 
mux_module mux_module_inst_1_2567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111])); 
fsm fsm_inst_1_2569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
fsm fsm_inst_1_2570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109])); 
mux_module mux_module_inst_1_2571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107])); 
fsm fsm_inst_1_2573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106])); 
mux_module mux_module_inst_1_2574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
fsm fsm_inst_1_2577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102])); 
mux_module mux_module_inst_1_2578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99])); 
fsm fsm_inst_1_2581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
mux_module mux_module_inst_1_2582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96])); 
mux_module mux_module_inst_1_2584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94])); 
mux_module mux_module_inst_1_2586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
fsm fsm_inst_1_2588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91])); 
fsm fsm_inst_1_2589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90])); 
mux_module mux_module_inst_1_2590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86])); 
fsm fsm_inst_1_2594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
mux_module mux_module_inst_1_2595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
mux_module mux_module_inst_1_2597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
mux_module mux_module_inst_1_2599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
fsm fsm_inst_1_2601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78])); 
mux_module mux_module_inst_1_2602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76])); 
fsm fsm_inst_1_2604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75])); 
fsm fsm_inst_1_2605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74])); 
mux_module mux_module_inst_1_2606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
mux_module mux_module_inst_1_2608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
fsm fsm_inst_1_2610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
mux_module mux_module_inst_1_2611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
fsm fsm_inst_1_2613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_2614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60])); 
mux_module mux_module_inst_1_2620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58])); 
mux_module mux_module_inst_1_2622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51])); 
fsm fsm_inst_1_2629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_2630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
mux_module mux_module_inst_1_2631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
mux_module mux_module_inst_1_2635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43])); 
fsm fsm_inst_1_2637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
fsm fsm_inst_1_2638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
mux_module mux_module_inst_1_2639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39])); 
mux_module mux_module_inst_1_2641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35])); 
fsm fsm_inst_1_2645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
mux_module mux_module_inst_1_2646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32])); 
mux_module mux_module_inst_1_2648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30])); 
mux_module mux_module_inst_1_2650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27])); 
fsm fsm_inst_1_2653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
fsm fsm_inst_1_2654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25])); 
fsm fsm_inst_1_2655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
fsm fsm_inst_1_2656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
mux_module mux_module_inst_1_2657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20])); 
mux_module mux_module_inst_1_2660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17])); 
fsm fsm_inst_1_2663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16])); 
mux_module mux_module_inst_1_2664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14])); 
mux_module mux_module_inst_1_2666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12])); 
fsm fsm_inst_1_2668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11])); 
fsm fsm_inst_1_2669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10])); 
mux_module mux_module_inst_1_2670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_2671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
fsm fsm_inst_1_2673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
fsm fsm_inst_1_2674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_2675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
mux_module mux_module_inst_1_2676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_2677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2])); 
fsm fsm_inst_1_2678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
mux_module mux_module_inst_1_2679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
always@(posedge clk) begin 
outp [2679:0] <= intermediate_reg_1; 
outp[4319:2680] <= intermediate_reg_1[1639:0] ; 
end 
endmodule 
 

module interface_27(input reg [3599:0] inp, output reg [1547:0] outp, input clk, input reset);
reg [3599:0]intermediate_reg_0; 
always@(posedge clk) begin 
intermediate_reg_0 <= inp; 
end 
 
reg [1799:0]intermediate_reg_1; 
 
mux_module mux_module_inst_1_0(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3599]),.i2(intermediate_reg_0[3598]),.o(intermediate_reg_1[1799]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3597]),.i2(intermediate_reg_0[3596]),.o(intermediate_reg_1[1798])); 
mux_module mux_module_inst_1_2(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3595]),.i2(intermediate_reg_0[3594]),.o(intermediate_reg_1[1797]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_3(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3593]),.i2(intermediate_reg_0[3592]),.o(intermediate_reg_1[1796]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_4(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3591]),.i2(intermediate_reg_0[3590]),.o(intermediate_reg_1[1795]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_5(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3589]),.i2(intermediate_reg_0[3588]),.o(intermediate_reg_1[1794]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_6(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3587]),.i2(intermediate_reg_0[3586]),.o(intermediate_reg_1[1793])); 
fsm fsm_inst_1_7(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3585]),.i2(intermediate_reg_0[3584]),.o(intermediate_reg_1[1792])); 
mux_module mux_module_inst_1_8(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3583]),.i2(intermediate_reg_0[3582]),.o(intermediate_reg_1[1791]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_9(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3581]),.i2(intermediate_reg_0[3580]),.o(intermediate_reg_1[1790])); 
mux_module mux_module_inst_1_10(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3579]),.i2(intermediate_reg_0[3578]),.o(intermediate_reg_1[1789]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_11(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3577]),.i2(intermediate_reg_0[3576]),.o(intermediate_reg_1[1788])); 
fsm fsm_inst_1_12(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3575]),.i2(intermediate_reg_0[3574]),.o(intermediate_reg_1[1787])); 
mux_module mux_module_inst_1_13(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3573]),.i2(intermediate_reg_0[3572]),.o(intermediate_reg_1[1786]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_14(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3571]),.i2(intermediate_reg_0[3570]),.o(intermediate_reg_1[1785]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_15(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3569]),.i2(intermediate_reg_0[3568]),.o(intermediate_reg_1[1784])); 
fsm fsm_inst_1_16(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3567]),.i2(intermediate_reg_0[3566]),.o(intermediate_reg_1[1783])); 
fsm fsm_inst_1_17(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3565]),.i2(intermediate_reg_0[3564]),.o(intermediate_reg_1[1782])); 
mux_module mux_module_inst_1_18(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3563]),.i2(intermediate_reg_0[3562]),.o(intermediate_reg_1[1781]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_19(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3561]),.i2(intermediate_reg_0[3560]),.o(intermediate_reg_1[1780])); 
fsm fsm_inst_1_20(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3559]),.i2(intermediate_reg_0[3558]),.o(intermediate_reg_1[1779])); 
fsm fsm_inst_1_21(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3557]),.i2(intermediate_reg_0[3556]),.o(intermediate_reg_1[1778])); 
mux_module mux_module_inst_1_22(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3555]),.i2(intermediate_reg_0[3554]),.o(intermediate_reg_1[1777]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_23(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3553]),.i2(intermediate_reg_0[3552]),.o(intermediate_reg_1[1776])); 
fsm fsm_inst_1_24(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3551]),.i2(intermediate_reg_0[3550]),.o(intermediate_reg_1[1775])); 
mux_module mux_module_inst_1_25(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3549]),.i2(intermediate_reg_0[3548]),.o(intermediate_reg_1[1774]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_26(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3547]),.i2(intermediate_reg_0[3546]),.o(intermediate_reg_1[1773])); 
mux_module mux_module_inst_1_27(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3545]),.i2(intermediate_reg_0[3544]),.o(intermediate_reg_1[1772]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_28(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3543]),.i2(intermediate_reg_0[3542]),.o(intermediate_reg_1[1771]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_29(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3541]),.i2(intermediate_reg_0[3540]),.o(intermediate_reg_1[1770]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_30(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3539]),.i2(intermediate_reg_0[3538]),.o(intermediate_reg_1[1769]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_31(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3537]),.i2(intermediate_reg_0[3536]),.o(intermediate_reg_1[1768])); 
fsm fsm_inst_1_32(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3535]),.i2(intermediate_reg_0[3534]),.o(intermediate_reg_1[1767])); 
mux_module mux_module_inst_1_33(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3533]),.i2(intermediate_reg_0[3532]),.o(intermediate_reg_1[1766]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_34(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3531]),.i2(intermediate_reg_0[3530]),.o(intermediate_reg_1[1765]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_35(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3529]),.i2(intermediate_reg_0[3528]),.o(intermediate_reg_1[1764])); 
mux_module mux_module_inst_1_36(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3527]),.i2(intermediate_reg_0[3526]),.o(intermediate_reg_1[1763]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_37(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3525]),.i2(intermediate_reg_0[3524]),.o(intermediate_reg_1[1762])); 
mux_module mux_module_inst_1_38(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3523]),.i2(intermediate_reg_0[3522]),.o(intermediate_reg_1[1761]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_39(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3521]),.i2(intermediate_reg_0[3520]),.o(intermediate_reg_1[1760]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_40(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3519]),.i2(intermediate_reg_0[3518]),.o(intermediate_reg_1[1759]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_41(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3517]),.i2(intermediate_reg_0[3516]),.o(intermediate_reg_1[1758])); 
mux_module mux_module_inst_1_42(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3515]),.i2(intermediate_reg_0[3514]),.o(intermediate_reg_1[1757]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_43(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3513]),.i2(intermediate_reg_0[3512]),.o(intermediate_reg_1[1756]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_44(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3511]),.i2(intermediate_reg_0[3510]),.o(intermediate_reg_1[1755]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_45(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3509]),.i2(intermediate_reg_0[3508]),.o(intermediate_reg_1[1754]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_46(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3507]),.i2(intermediate_reg_0[3506]),.o(intermediate_reg_1[1753]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_47(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3505]),.i2(intermediate_reg_0[3504]),.o(intermediate_reg_1[1752]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_48(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3503]),.i2(intermediate_reg_0[3502]),.o(intermediate_reg_1[1751])); 
fsm fsm_inst_1_49(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3501]),.i2(intermediate_reg_0[3500]),.o(intermediate_reg_1[1750])); 
mux_module mux_module_inst_1_50(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3499]),.i2(intermediate_reg_0[3498]),.o(intermediate_reg_1[1749]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_51(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3497]),.i2(intermediate_reg_0[3496]),.o(intermediate_reg_1[1748]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_52(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3495]),.i2(intermediate_reg_0[3494]),.o(intermediate_reg_1[1747])); 
fsm fsm_inst_1_53(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3493]),.i2(intermediate_reg_0[3492]),.o(intermediate_reg_1[1746])); 
mux_module mux_module_inst_1_54(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3491]),.i2(intermediate_reg_0[3490]),.o(intermediate_reg_1[1745]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_55(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3489]),.i2(intermediate_reg_0[3488]),.o(intermediate_reg_1[1744]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_56(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3487]),.i2(intermediate_reg_0[3486]),.o(intermediate_reg_1[1743])); 
fsm fsm_inst_1_57(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3485]),.i2(intermediate_reg_0[3484]),.o(intermediate_reg_1[1742])); 
mux_module mux_module_inst_1_58(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3483]),.i2(intermediate_reg_0[3482]),.o(intermediate_reg_1[1741]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_59(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3481]),.i2(intermediate_reg_0[3480]),.o(intermediate_reg_1[1740]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_60(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3479]),.i2(intermediate_reg_0[3478]),.o(intermediate_reg_1[1739])); 
fsm fsm_inst_1_61(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3477]),.i2(intermediate_reg_0[3476]),.o(intermediate_reg_1[1738])); 
fsm fsm_inst_1_62(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3475]),.i2(intermediate_reg_0[3474]),.o(intermediate_reg_1[1737])); 
fsm fsm_inst_1_63(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3473]),.i2(intermediate_reg_0[3472]),.o(intermediate_reg_1[1736])); 
mux_module mux_module_inst_1_64(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3471]),.i2(intermediate_reg_0[3470]),.o(intermediate_reg_1[1735]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_65(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3469]),.i2(intermediate_reg_0[3468]),.o(intermediate_reg_1[1734])); 
fsm fsm_inst_1_66(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3467]),.i2(intermediate_reg_0[3466]),.o(intermediate_reg_1[1733])); 
mux_module mux_module_inst_1_67(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3465]),.i2(intermediate_reg_0[3464]),.o(intermediate_reg_1[1732]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_68(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3463]),.i2(intermediate_reg_0[3462]),.o(intermediate_reg_1[1731])); 
fsm fsm_inst_1_69(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3461]),.i2(intermediate_reg_0[3460]),.o(intermediate_reg_1[1730])); 
mux_module mux_module_inst_1_70(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3459]),.i2(intermediate_reg_0[3458]),.o(intermediate_reg_1[1729]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_71(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3457]),.i2(intermediate_reg_0[3456]),.o(intermediate_reg_1[1728]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_72(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3455]),.i2(intermediate_reg_0[3454]),.o(intermediate_reg_1[1727])); 
mux_module mux_module_inst_1_73(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3453]),.i2(intermediate_reg_0[3452]),.o(intermediate_reg_1[1726]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_74(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3451]),.i2(intermediate_reg_0[3450]),.o(intermediate_reg_1[1725]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_75(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3449]),.i2(intermediate_reg_0[3448]),.o(intermediate_reg_1[1724]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_76(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3447]),.i2(intermediate_reg_0[3446]),.o(intermediate_reg_1[1723]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_77(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3445]),.i2(intermediate_reg_0[3444]),.o(intermediate_reg_1[1722])); 
mux_module mux_module_inst_1_78(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3443]),.i2(intermediate_reg_0[3442]),.o(intermediate_reg_1[1721]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_79(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3441]),.i2(intermediate_reg_0[3440]),.o(intermediate_reg_1[1720])); 
fsm fsm_inst_1_80(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3439]),.i2(intermediate_reg_0[3438]),.o(intermediate_reg_1[1719])); 
mux_module mux_module_inst_1_81(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3437]),.i2(intermediate_reg_0[3436]),.o(intermediate_reg_1[1718]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_82(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3435]),.i2(intermediate_reg_0[3434]),.o(intermediate_reg_1[1717]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_83(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3433]),.i2(intermediate_reg_0[3432]),.o(intermediate_reg_1[1716]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_84(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3431]),.i2(intermediate_reg_0[3430]),.o(intermediate_reg_1[1715]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_85(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3429]),.i2(intermediate_reg_0[3428]),.o(intermediate_reg_1[1714]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_86(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3427]),.i2(intermediate_reg_0[3426]),.o(intermediate_reg_1[1713])); 
fsm fsm_inst_1_87(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3425]),.i2(intermediate_reg_0[3424]),.o(intermediate_reg_1[1712])); 
fsm fsm_inst_1_88(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3423]),.i2(intermediate_reg_0[3422]),.o(intermediate_reg_1[1711])); 
fsm fsm_inst_1_89(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3421]),.i2(intermediate_reg_0[3420]),.o(intermediate_reg_1[1710])); 
fsm fsm_inst_1_90(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3419]),.i2(intermediate_reg_0[3418]),.o(intermediate_reg_1[1709])); 
fsm fsm_inst_1_91(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3417]),.i2(intermediate_reg_0[3416]),.o(intermediate_reg_1[1708])); 
mux_module mux_module_inst_1_92(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3415]),.i2(intermediate_reg_0[3414]),.o(intermediate_reg_1[1707]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_93(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3413]),.i2(intermediate_reg_0[3412]),.o(intermediate_reg_1[1706]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_94(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3411]),.i2(intermediate_reg_0[3410]),.o(intermediate_reg_1[1705]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_95(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3409]),.i2(intermediate_reg_0[3408]),.o(intermediate_reg_1[1704]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_96(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3407]),.i2(intermediate_reg_0[3406]),.o(intermediate_reg_1[1703])); 
fsm fsm_inst_1_97(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3405]),.i2(intermediate_reg_0[3404]),.o(intermediate_reg_1[1702])); 
mux_module mux_module_inst_1_98(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3403]),.i2(intermediate_reg_0[3402]),.o(intermediate_reg_1[1701]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_99(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3401]),.i2(intermediate_reg_0[3400]),.o(intermediate_reg_1[1700])); 
fsm fsm_inst_1_100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3399]),.i2(intermediate_reg_0[3398]),.o(intermediate_reg_1[1699])); 
mux_module mux_module_inst_1_101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3397]),.i2(intermediate_reg_0[3396]),.o(intermediate_reg_1[1698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3395]),.i2(intermediate_reg_0[3394]),.o(intermediate_reg_1[1697]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3393]),.i2(intermediate_reg_0[3392]),.o(intermediate_reg_1[1696]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3391]),.i2(intermediate_reg_0[3390]),.o(intermediate_reg_1[1695])); 
fsm fsm_inst_1_105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3389]),.i2(intermediate_reg_0[3388]),.o(intermediate_reg_1[1694])); 
fsm fsm_inst_1_106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3387]),.i2(intermediate_reg_0[3386]),.o(intermediate_reg_1[1693])); 
mux_module mux_module_inst_1_107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3385]),.i2(intermediate_reg_0[3384]),.o(intermediate_reg_1[1692]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3383]),.i2(intermediate_reg_0[3382]),.o(intermediate_reg_1[1691]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3381]),.i2(intermediate_reg_0[3380]),.o(intermediate_reg_1[1690]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3379]),.i2(intermediate_reg_0[3378]),.o(intermediate_reg_1[1689]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3377]),.i2(intermediate_reg_0[3376]),.o(intermediate_reg_1[1688]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3375]),.i2(intermediate_reg_0[3374]),.o(intermediate_reg_1[1687])); 
mux_module mux_module_inst_1_113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3373]),.i2(intermediate_reg_0[3372]),.o(intermediate_reg_1[1686]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3371]),.i2(intermediate_reg_0[3370]),.o(intermediate_reg_1[1685]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3369]),.i2(intermediate_reg_0[3368]),.o(intermediate_reg_1[1684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3367]),.i2(intermediate_reg_0[3366]),.o(intermediate_reg_1[1683]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3365]),.i2(intermediate_reg_0[3364]),.o(intermediate_reg_1[1682])); 
fsm fsm_inst_1_118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3363]),.i2(intermediate_reg_0[3362]),.o(intermediate_reg_1[1681])); 
mux_module mux_module_inst_1_119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3361]),.i2(intermediate_reg_0[3360]),.o(intermediate_reg_1[1680]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3359]),.i2(intermediate_reg_0[3358]),.o(intermediate_reg_1[1679]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3357]),.i2(intermediate_reg_0[3356]),.o(intermediate_reg_1[1678])); 
fsm fsm_inst_1_122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3355]),.i2(intermediate_reg_0[3354]),.o(intermediate_reg_1[1677])); 
fsm fsm_inst_1_123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3353]),.i2(intermediate_reg_0[3352]),.o(intermediate_reg_1[1676])); 
mux_module mux_module_inst_1_124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3351]),.i2(intermediate_reg_0[3350]),.o(intermediate_reg_1[1675]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3349]),.i2(intermediate_reg_0[3348]),.o(intermediate_reg_1[1674]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3347]),.i2(intermediate_reg_0[3346]),.o(intermediate_reg_1[1673]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3345]),.i2(intermediate_reg_0[3344]),.o(intermediate_reg_1[1672]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3343]),.i2(intermediate_reg_0[3342]),.o(intermediate_reg_1[1671]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3341]),.i2(intermediate_reg_0[3340]),.o(intermediate_reg_1[1670]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3339]),.i2(intermediate_reg_0[3338]),.o(intermediate_reg_1[1669]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3337]),.i2(intermediate_reg_0[3336]),.o(intermediate_reg_1[1668])); 
mux_module mux_module_inst_1_132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3335]),.i2(intermediate_reg_0[3334]),.o(intermediate_reg_1[1667]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3333]),.i2(intermediate_reg_0[3332]),.o(intermediate_reg_1[1666])); 
mux_module mux_module_inst_1_134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3331]),.i2(intermediate_reg_0[3330]),.o(intermediate_reg_1[1665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3329]),.i2(intermediate_reg_0[3328]),.o(intermediate_reg_1[1664]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3327]),.i2(intermediate_reg_0[3326]),.o(intermediate_reg_1[1663])); 
mux_module mux_module_inst_1_137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3325]),.i2(intermediate_reg_0[3324]),.o(intermediate_reg_1[1662]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3323]),.i2(intermediate_reg_0[3322]),.o(intermediate_reg_1[1661]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3321]),.i2(intermediate_reg_0[3320]),.o(intermediate_reg_1[1660])); 
fsm fsm_inst_1_140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3319]),.i2(intermediate_reg_0[3318]),.o(intermediate_reg_1[1659])); 
fsm fsm_inst_1_141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3317]),.i2(intermediate_reg_0[3316]),.o(intermediate_reg_1[1658])); 
fsm fsm_inst_1_142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3315]),.i2(intermediate_reg_0[3314]),.o(intermediate_reg_1[1657])); 
fsm fsm_inst_1_143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3313]),.i2(intermediate_reg_0[3312]),.o(intermediate_reg_1[1656])); 
mux_module mux_module_inst_1_144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3311]),.i2(intermediate_reg_0[3310]),.o(intermediate_reg_1[1655]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3309]),.i2(intermediate_reg_0[3308]),.o(intermediate_reg_1[1654]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3307]),.i2(intermediate_reg_0[3306]),.o(intermediate_reg_1[1653])); 
fsm fsm_inst_1_147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3305]),.i2(intermediate_reg_0[3304]),.o(intermediate_reg_1[1652])); 
fsm fsm_inst_1_148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3303]),.i2(intermediate_reg_0[3302]),.o(intermediate_reg_1[1651])); 
fsm fsm_inst_1_149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3301]),.i2(intermediate_reg_0[3300]),.o(intermediate_reg_1[1650])); 
mux_module mux_module_inst_1_150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3299]),.i2(intermediate_reg_0[3298]),.o(intermediate_reg_1[1649]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3297]),.i2(intermediate_reg_0[3296]),.o(intermediate_reg_1[1648])); 
fsm fsm_inst_1_152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3295]),.i2(intermediate_reg_0[3294]),.o(intermediate_reg_1[1647])); 
fsm fsm_inst_1_153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3293]),.i2(intermediate_reg_0[3292]),.o(intermediate_reg_1[1646])); 
fsm fsm_inst_1_154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3291]),.i2(intermediate_reg_0[3290]),.o(intermediate_reg_1[1645])); 
fsm fsm_inst_1_155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3289]),.i2(intermediate_reg_0[3288]),.o(intermediate_reg_1[1644])); 
mux_module mux_module_inst_1_156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3287]),.i2(intermediate_reg_0[3286]),.o(intermediate_reg_1[1643]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3285]),.i2(intermediate_reg_0[3284]),.o(intermediate_reg_1[1642]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3283]),.i2(intermediate_reg_0[3282]),.o(intermediate_reg_1[1641])); 
fsm fsm_inst_1_159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3281]),.i2(intermediate_reg_0[3280]),.o(intermediate_reg_1[1640])); 
fsm fsm_inst_1_160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3279]),.i2(intermediate_reg_0[3278]),.o(intermediate_reg_1[1639])); 
fsm fsm_inst_1_161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3277]),.i2(intermediate_reg_0[3276]),.o(intermediate_reg_1[1638])); 
mux_module mux_module_inst_1_162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3275]),.i2(intermediate_reg_0[3274]),.o(intermediate_reg_1[1637]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3273]),.i2(intermediate_reg_0[3272]),.o(intermediate_reg_1[1636])); 
fsm fsm_inst_1_164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3271]),.i2(intermediate_reg_0[3270]),.o(intermediate_reg_1[1635])); 
mux_module mux_module_inst_1_165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3269]),.i2(intermediate_reg_0[3268]),.o(intermediate_reg_1[1634]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3267]),.i2(intermediate_reg_0[3266]),.o(intermediate_reg_1[1633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3265]),.i2(intermediate_reg_0[3264]),.o(intermediate_reg_1[1632]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3263]),.i2(intermediate_reg_0[3262]),.o(intermediate_reg_1[1631]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3261]),.i2(intermediate_reg_0[3260]),.o(intermediate_reg_1[1630]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3259]),.i2(intermediate_reg_0[3258]),.o(intermediate_reg_1[1629])); 
mux_module mux_module_inst_1_171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3257]),.i2(intermediate_reg_0[3256]),.o(intermediate_reg_1[1628]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3255]),.i2(intermediate_reg_0[3254]),.o(intermediate_reg_1[1627])); 
fsm fsm_inst_1_173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3253]),.i2(intermediate_reg_0[3252]),.o(intermediate_reg_1[1626])); 
mux_module mux_module_inst_1_174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3251]),.i2(intermediate_reg_0[3250]),.o(intermediate_reg_1[1625]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3249]),.i2(intermediate_reg_0[3248]),.o(intermediate_reg_1[1624])); 
fsm fsm_inst_1_176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3247]),.i2(intermediate_reg_0[3246]),.o(intermediate_reg_1[1623])); 
mux_module mux_module_inst_1_177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3245]),.i2(intermediate_reg_0[3244]),.o(intermediate_reg_1[1622]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3243]),.i2(intermediate_reg_0[3242]),.o(intermediate_reg_1[1621])); 
mux_module mux_module_inst_1_179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3241]),.i2(intermediate_reg_0[3240]),.o(intermediate_reg_1[1620]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3239]),.i2(intermediate_reg_0[3238]),.o(intermediate_reg_1[1619]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3237]),.i2(intermediate_reg_0[3236]),.o(intermediate_reg_1[1618]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3235]),.i2(intermediate_reg_0[3234]),.o(intermediate_reg_1[1617]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3233]),.i2(intermediate_reg_0[3232]),.o(intermediate_reg_1[1616]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3231]),.i2(intermediate_reg_0[3230]),.o(intermediate_reg_1[1615])); 
mux_module mux_module_inst_1_185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3229]),.i2(intermediate_reg_0[3228]),.o(intermediate_reg_1[1614]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3227]),.i2(intermediate_reg_0[3226]),.o(intermediate_reg_1[1613]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3225]),.i2(intermediate_reg_0[3224]),.o(intermediate_reg_1[1612])); 
mux_module mux_module_inst_1_188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3223]),.i2(intermediate_reg_0[3222]),.o(intermediate_reg_1[1611]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3221]),.i2(intermediate_reg_0[3220]),.o(intermediate_reg_1[1610])); 
fsm fsm_inst_1_190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3219]),.i2(intermediate_reg_0[3218]),.o(intermediate_reg_1[1609])); 
fsm fsm_inst_1_191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3217]),.i2(intermediate_reg_0[3216]),.o(intermediate_reg_1[1608])); 
mux_module mux_module_inst_1_192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3215]),.i2(intermediate_reg_0[3214]),.o(intermediate_reg_1[1607]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3213]),.i2(intermediate_reg_0[3212]),.o(intermediate_reg_1[1606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3211]),.i2(intermediate_reg_0[3210]),.o(intermediate_reg_1[1605]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3209]),.i2(intermediate_reg_0[3208]),.o(intermediate_reg_1[1604])); 
fsm fsm_inst_1_196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3207]),.i2(intermediate_reg_0[3206]),.o(intermediate_reg_1[1603])); 
mux_module mux_module_inst_1_197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3205]),.i2(intermediate_reg_0[3204]),.o(intermediate_reg_1[1602]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3203]),.i2(intermediate_reg_0[3202]),.o(intermediate_reg_1[1601]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3201]),.i2(intermediate_reg_0[3200]),.o(intermediate_reg_1[1600]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3199]),.i2(intermediate_reg_0[3198]),.o(intermediate_reg_1[1599])); 
fsm fsm_inst_1_201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3197]),.i2(intermediate_reg_0[3196]),.o(intermediate_reg_1[1598])); 
mux_module mux_module_inst_1_202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3195]),.i2(intermediate_reg_0[3194]),.o(intermediate_reg_1[1597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3193]),.i2(intermediate_reg_0[3192]),.o(intermediate_reg_1[1596]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3191]),.i2(intermediate_reg_0[3190]),.o(intermediate_reg_1[1595]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3189]),.i2(intermediate_reg_0[3188]),.o(intermediate_reg_1[1594])); 
mux_module mux_module_inst_1_206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3187]),.i2(intermediate_reg_0[3186]),.o(intermediate_reg_1[1593]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3185]),.i2(intermediate_reg_0[3184]),.o(intermediate_reg_1[1592]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3183]),.i2(intermediate_reg_0[3182]),.o(intermediate_reg_1[1591])); 
fsm fsm_inst_1_209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3181]),.i2(intermediate_reg_0[3180]),.o(intermediate_reg_1[1590])); 
mux_module mux_module_inst_1_210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3179]),.i2(intermediate_reg_0[3178]),.o(intermediate_reg_1[1589]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3177]),.i2(intermediate_reg_0[3176]),.o(intermediate_reg_1[1588])); 
mux_module mux_module_inst_1_212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3175]),.i2(intermediate_reg_0[3174]),.o(intermediate_reg_1[1587]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3173]),.i2(intermediate_reg_0[3172]),.o(intermediate_reg_1[1586]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3171]),.i2(intermediate_reg_0[3170]),.o(intermediate_reg_1[1585]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3169]),.i2(intermediate_reg_0[3168]),.o(intermediate_reg_1[1584]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3167]),.i2(intermediate_reg_0[3166]),.o(intermediate_reg_1[1583]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3165]),.i2(intermediate_reg_0[3164]),.o(intermediate_reg_1[1582]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3163]),.i2(intermediate_reg_0[3162]),.o(intermediate_reg_1[1581])); 
fsm fsm_inst_1_219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3161]),.i2(intermediate_reg_0[3160]),.o(intermediate_reg_1[1580])); 
mux_module mux_module_inst_1_220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3159]),.i2(intermediate_reg_0[3158]),.o(intermediate_reg_1[1579]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3157]),.i2(intermediate_reg_0[3156]),.o(intermediate_reg_1[1578]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3155]),.i2(intermediate_reg_0[3154]),.o(intermediate_reg_1[1577]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3153]),.i2(intermediate_reg_0[3152]),.o(intermediate_reg_1[1576]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3151]),.i2(intermediate_reg_0[3150]),.o(intermediate_reg_1[1575])); 
fsm fsm_inst_1_225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3149]),.i2(intermediate_reg_0[3148]),.o(intermediate_reg_1[1574])); 
mux_module mux_module_inst_1_226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3147]),.i2(intermediate_reg_0[3146]),.o(intermediate_reg_1[1573]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3145]),.i2(intermediate_reg_0[3144]),.o(intermediate_reg_1[1572])); 
mux_module mux_module_inst_1_228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3143]),.i2(intermediate_reg_0[3142]),.o(intermediate_reg_1[1571]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3141]),.i2(intermediate_reg_0[3140]),.o(intermediate_reg_1[1570]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3139]),.i2(intermediate_reg_0[3138]),.o(intermediate_reg_1[1569])); 
fsm fsm_inst_1_231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3137]),.i2(intermediate_reg_0[3136]),.o(intermediate_reg_1[1568])); 
mux_module mux_module_inst_1_232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3135]),.i2(intermediate_reg_0[3134]),.o(intermediate_reg_1[1567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3133]),.i2(intermediate_reg_0[3132]),.o(intermediate_reg_1[1566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3131]),.i2(intermediate_reg_0[3130]),.o(intermediate_reg_1[1565]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3129]),.i2(intermediate_reg_0[3128]),.o(intermediate_reg_1[1564])); 
fsm fsm_inst_1_236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3127]),.i2(intermediate_reg_0[3126]),.o(intermediate_reg_1[1563])); 
fsm fsm_inst_1_237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3125]),.i2(intermediate_reg_0[3124]),.o(intermediate_reg_1[1562])); 
mux_module mux_module_inst_1_238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3123]),.i2(intermediate_reg_0[3122]),.o(intermediate_reg_1[1561]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3121]),.i2(intermediate_reg_0[3120]),.o(intermediate_reg_1[1560])); 
fsm fsm_inst_1_240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3119]),.i2(intermediate_reg_0[3118]),.o(intermediate_reg_1[1559])); 
fsm fsm_inst_1_241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3117]),.i2(intermediate_reg_0[3116]),.o(intermediate_reg_1[1558])); 
fsm fsm_inst_1_242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3115]),.i2(intermediate_reg_0[3114]),.o(intermediate_reg_1[1557])); 
mux_module mux_module_inst_1_243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3113]),.i2(intermediate_reg_0[3112]),.o(intermediate_reg_1[1556]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3111]),.i2(intermediate_reg_0[3110]),.o(intermediate_reg_1[1555]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3109]),.i2(intermediate_reg_0[3108]),.o(intermediate_reg_1[1554])); 
mux_module mux_module_inst_1_246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3107]),.i2(intermediate_reg_0[3106]),.o(intermediate_reg_1[1553]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3105]),.i2(intermediate_reg_0[3104]),.o(intermediate_reg_1[1552]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3103]),.i2(intermediate_reg_0[3102]),.o(intermediate_reg_1[1551]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3101]),.i2(intermediate_reg_0[3100]),.o(intermediate_reg_1[1550])); 
mux_module mux_module_inst_1_250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3099]),.i2(intermediate_reg_0[3098]),.o(intermediate_reg_1[1549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3097]),.i2(intermediate_reg_0[3096]),.o(intermediate_reg_1[1548]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3095]),.i2(intermediate_reg_0[3094]),.o(intermediate_reg_1[1547])); 
fsm fsm_inst_1_253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3093]),.i2(intermediate_reg_0[3092]),.o(intermediate_reg_1[1546])); 
fsm fsm_inst_1_254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3091]),.i2(intermediate_reg_0[3090]),.o(intermediate_reg_1[1545])); 
mux_module mux_module_inst_1_255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3089]),.i2(intermediate_reg_0[3088]),.o(intermediate_reg_1[1544]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3087]),.i2(intermediate_reg_0[3086]),.o(intermediate_reg_1[1543])); 
mux_module mux_module_inst_1_257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3085]),.i2(intermediate_reg_0[3084]),.o(intermediate_reg_1[1542]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3083]),.i2(intermediate_reg_0[3082]),.o(intermediate_reg_1[1541]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3081]),.i2(intermediate_reg_0[3080]),.o(intermediate_reg_1[1540]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3079]),.i2(intermediate_reg_0[3078]),.o(intermediate_reg_1[1539]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3077]),.i2(intermediate_reg_0[3076]),.o(intermediate_reg_1[1538])); 
fsm fsm_inst_1_262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3075]),.i2(intermediate_reg_0[3074]),.o(intermediate_reg_1[1537])); 
fsm fsm_inst_1_263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3073]),.i2(intermediate_reg_0[3072]),.o(intermediate_reg_1[1536])); 
fsm fsm_inst_1_264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3071]),.i2(intermediate_reg_0[3070]),.o(intermediate_reg_1[1535])); 
mux_module mux_module_inst_1_265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3069]),.i2(intermediate_reg_0[3068]),.o(intermediate_reg_1[1534]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3067]),.i2(intermediate_reg_0[3066]),.o(intermediate_reg_1[1533])); 
mux_module mux_module_inst_1_267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3065]),.i2(intermediate_reg_0[3064]),.o(intermediate_reg_1[1532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3063]),.i2(intermediate_reg_0[3062]),.o(intermediate_reg_1[1531]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3061]),.i2(intermediate_reg_0[3060]),.o(intermediate_reg_1[1530])); 
mux_module mux_module_inst_1_270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3059]),.i2(intermediate_reg_0[3058]),.o(intermediate_reg_1[1529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3057]),.i2(intermediate_reg_0[3056]),.o(intermediate_reg_1[1528]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3055]),.i2(intermediate_reg_0[3054]),.o(intermediate_reg_1[1527])); 
mux_module mux_module_inst_1_273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3053]),.i2(intermediate_reg_0[3052]),.o(intermediate_reg_1[1526]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3051]),.i2(intermediate_reg_0[3050]),.o(intermediate_reg_1[1525])); 
mux_module mux_module_inst_1_275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3049]),.i2(intermediate_reg_0[3048]),.o(intermediate_reg_1[1524]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3047]),.i2(intermediate_reg_0[3046]),.o(intermediate_reg_1[1523])); 
fsm fsm_inst_1_277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3045]),.i2(intermediate_reg_0[3044]),.o(intermediate_reg_1[1522])); 
fsm fsm_inst_1_278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3043]),.i2(intermediate_reg_0[3042]),.o(intermediate_reg_1[1521])); 
fsm fsm_inst_1_279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3041]),.i2(intermediate_reg_0[3040]),.o(intermediate_reg_1[1520])); 
mux_module mux_module_inst_1_280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3039]),.i2(intermediate_reg_0[3038]),.o(intermediate_reg_1[1519]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3037]),.i2(intermediate_reg_0[3036]),.o(intermediate_reg_1[1518]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3035]),.i2(intermediate_reg_0[3034]),.o(intermediate_reg_1[1517])); 
fsm fsm_inst_1_283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3033]),.i2(intermediate_reg_0[3032]),.o(intermediate_reg_1[1516])); 
fsm fsm_inst_1_284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3031]),.i2(intermediate_reg_0[3030]),.o(intermediate_reg_1[1515])); 
fsm fsm_inst_1_285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3029]),.i2(intermediate_reg_0[3028]),.o(intermediate_reg_1[1514])); 
mux_module mux_module_inst_1_286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3027]),.i2(intermediate_reg_0[3026]),.o(intermediate_reg_1[1513]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3025]),.i2(intermediate_reg_0[3024]),.o(intermediate_reg_1[1512]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3023]),.i2(intermediate_reg_0[3022]),.o(intermediate_reg_1[1511])); 
fsm fsm_inst_1_289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3021]),.i2(intermediate_reg_0[3020]),.o(intermediate_reg_1[1510])); 
mux_module mux_module_inst_1_290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3019]),.i2(intermediate_reg_0[3018]),.o(intermediate_reg_1[1509]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3017]),.i2(intermediate_reg_0[3016]),.o(intermediate_reg_1[1508])); 
fsm fsm_inst_1_292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3015]),.i2(intermediate_reg_0[3014]),.o(intermediate_reg_1[1507])); 
fsm fsm_inst_1_293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3013]),.i2(intermediate_reg_0[3012]),.o(intermediate_reg_1[1506])); 
fsm fsm_inst_1_294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3011]),.i2(intermediate_reg_0[3010]),.o(intermediate_reg_1[1505])); 
mux_module mux_module_inst_1_295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3009]),.i2(intermediate_reg_0[3008]),.o(intermediate_reg_1[1504]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3007]),.i2(intermediate_reg_0[3006]),.o(intermediate_reg_1[1503])); 
fsm fsm_inst_1_297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3005]),.i2(intermediate_reg_0[3004]),.o(intermediate_reg_1[1502])); 
mux_module mux_module_inst_1_298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3003]),.i2(intermediate_reg_0[3002]),.o(intermediate_reg_1[1501]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3001]),.i2(intermediate_reg_0[3000]),.o(intermediate_reg_1[1500]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2999]),.i2(intermediate_reg_0[2998]),.o(intermediate_reg_1[1499])); 
mux_module mux_module_inst_1_301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2997]),.i2(intermediate_reg_0[2996]),.o(intermediate_reg_1[1498]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2995]),.i2(intermediate_reg_0[2994]),.o(intermediate_reg_1[1497])); 
mux_module mux_module_inst_1_303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2993]),.i2(intermediate_reg_0[2992]),.o(intermediate_reg_1[1496]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2991]),.i2(intermediate_reg_0[2990]),.o(intermediate_reg_1[1495]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2989]),.i2(intermediate_reg_0[2988]),.o(intermediate_reg_1[1494])); 
fsm fsm_inst_1_306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2987]),.i2(intermediate_reg_0[2986]),.o(intermediate_reg_1[1493])); 
fsm fsm_inst_1_307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2985]),.i2(intermediate_reg_0[2984]),.o(intermediate_reg_1[1492])); 
fsm fsm_inst_1_308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2983]),.i2(intermediate_reg_0[2982]),.o(intermediate_reg_1[1491])); 
fsm fsm_inst_1_309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2981]),.i2(intermediate_reg_0[2980]),.o(intermediate_reg_1[1490])); 
fsm fsm_inst_1_310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2979]),.i2(intermediate_reg_0[2978]),.o(intermediate_reg_1[1489])); 
fsm fsm_inst_1_311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2977]),.i2(intermediate_reg_0[2976]),.o(intermediate_reg_1[1488])); 
mux_module mux_module_inst_1_312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2975]),.i2(intermediate_reg_0[2974]),.o(intermediate_reg_1[1487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2973]),.i2(intermediate_reg_0[2972]),.o(intermediate_reg_1[1486]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2971]),.i2(intermediate_reg_0[2970]),.o(intermediate_reg_1[1485]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2969]),.i2(intermediate_reg_0[2968]),.o(intermediate_reg_1[1484])); 
fsm fsm_inst_1_316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2967]),.i2(intermediate_reg_0[2966]),.o(intermediate_reg_1[1483])); 
mux_module mux_module_inst_1_317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2965]),.i2(intermediate_reg_0[2964]),.o(intermediate_reg_1[1482]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2963]),.i2(intermediate_reg_0[2962]),.o(intermediate_reg_1[1481]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2961]),.i2(intermediate_reg_0[2960]),.o(intermediate_reg_1[1480])); 
mux_module mux_module_inst_1_320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2959]),.i2(intermediate_reg_0[2958]),.o(intermediate_reg_1[1479]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2957]),.i2(intermediate_reg_0[2956]),.o(intermediate_reg_1[1478]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2955]),.i2(intermediate_reg_0[2954]),.o(intermediate_reg_1[1477]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2953]),.i2(intermediate_reg_0[2952]),.o(intermediate_reg_1[1476]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2951]),.i2(intermediate_reg_0[2950]),.o(intermediate_reg_1[1475])); 
fsm fsm_inst_1_325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2949]),.i2(intermediate_reg_0[2948]),.o(intermediate_reg_1[1474])); 
mux_module mux_module_inst_1_326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2947]),.i2(intermediate_reg_0[2946]),.o(intermediate_reg_1[1473]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2945]),.i2(intermediate_reg_0[2944]),.o(intermediate_reg_1[1472])); 
mux_module mux_module_inst_1_328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2943]),.i2(intermediate_reg_0[2942]),.o(intermediate_reg_1[1471]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2941]),.i2(intermediate_reg_0[2940]),.o(intermediate_reg_1[1470]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2939]),.i2(intermediate_reg_0[2938]),.o(intermediate_reg_1[1469]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2937]),.i2(intermediate_reg_0[2936]),.o(intermediate_reg_1[1468]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2935]),.i2(intermediate_reg_0[2934]),.o(intermediate_reg_1[1467]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2933]),.i2(intermediate_reg_0[2932]),.o(intermediate_reg_1[1466]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2931]),.i2(intermediate_reg_0[2930]),.o(intermediate_reg_1[1465]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2929]),.i2(intermediate_reg_0[2928]),.o(intermediate_reg_1[1464])); 
fsm fsm_inst_1_336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2927]),.i2(intermediate_reg_0[2926]),.o(intermediate_reg_1[1463])); 
fsm fsm_inst_1_337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2925]),.i2(intermediate_reg_0[2924]),.o(intermediate_reg_1[1462])); 
mux_module mux_module_inst_1_338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2923]),.i2(intermediate_reg_0[2922]),.o(intermediate_reg_1[1461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2921]),.i2(intermediate_reg_0[2920]),.o(intermediate_reg_1[1460]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2919]),.i2(intermediate_reg_0[2918]),.o(intermediate_reg_1[1459]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2917]),.i2(intermediate_reg_0[2916]),.o(intermediate_reg_1[1458]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2915]),.i2(intermediate_reg_0[2914]),.o(intermediate_reg_1[1457])); 
mux_module mux_module_inst_1_343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2913]),.i2(intermediate_reg_0[2912]),.o(intermediate_reg_1[1456]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2911]),.i2(intermediate_reg_0[2910]),.o(intermediate_reg_1[1455])); 
fsm fsm_inst_1_345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2909]),.i2(intermediate_reg_0[2908]),.o(intermediate_reg_1[1454])); 
mux_module mux_module_inst_1_346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2907]),.i2(intermediate_reg_0[2906]),.o(intermediate_reg_1[1453]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2905]),.i2(intermediate_reg_0[2904]),.o(intermediate_reg_1[1452]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2903]),.i2(intermediate_reg_0[2902]),.o(intermediate_reg_1[1451])); 
fsm fsm_inst_1_349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2901]),.i2(intermediate_reg_0[2900]),.o(intermediate_reg_1[1450])); 
fsm fsm_inst_1_350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2899]),.i2(intermediate_reg_0[2898]),.o(intermediate_reg_1[1449])); 
mux_module mux_module_inst_1_351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2897]),.i2(intermediate_reg_0[2896]),.o(intermediate_reg_1[1448]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2895]),.i2(intermediate_reg_0[2894]),.o(intermediate_reg_1[1447]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2893]),.i2(intermediate_reg_0[2892]),.o(intermediate_reg_1[1446])); 
fsm fsm_inst_1_354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2891]),.i2(intermediate_reg_0[2890]),.o(intermediate_reg_1[1445])); 
fsm fsm_inst_1_355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2889]),.i2(intermediate_reg_0[2888]),.o(intermediate_reg_1[1444])); 
fsm fsm_inst_1_356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2887]),.i2(intermediate_reg_0[2886]),.o(intermediate_reg_1[1443])); 
mux_module mux_module_inst_1_357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2885]),.i2(intermediate_reg_0[2884]),.o(intermediate_reg_1[1442]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2883]),.i2(intermediate_reg_0[2882]),.o(intermediate_reg_1[1441])); 
mux_module mux_module_inst_1_359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2881]),.i2(intermediate_reg_0[2880]),.o(intermediate_reg_1[1440]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2879]),.i2(intermediate_reg_0[2878]),.o(intermediate_reg_1[1439]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2877]),.i2(intermediate_reg_0[2876]),.o(intermediate_reg_1[1438])); 
fsm fsm_inst_1_362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2875]),.i2(intermediate_reg_0[2874]),.o(intermediate_reg_1[1437])); 
fsm fsm_inst_1_363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2873]),.i2(intermediate_reg_0[2872]),.o(intermediate_reg_1[1436])); 
fsm fsm_inst_1_364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2871]),.i2(intermediate_reg_0[2870]),.o(intermediate_reg_1[1435])); 
mux_module mux_module_inst_1_365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2869]),.i2(intermediate_reg_0[2868]),.o(intermediate_reg_1[1434]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2867]),.i2(intermediate_reg_0[2866]),.o(intermediate_reg_1[1433])); 
mux_module mux_module_inst_1_367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2865]),.i2(intermediate_reg_0[2864]),.o(intermediate_reg_1[1432]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2863]),.i2(intermediate_reg_0[2862]),.o(intermediate_reg_1[1431])); 
mux_module mux_module_inst_1_369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2861]),.i2(intermediate_reg_0[2860]),.o(intermediate_reg_1[1430]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2859]),.i2(intermediate_reg_0[2858]),.o(intermediate_reg_1[1429])); 
fsm fsm_inst_1_371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2857]),.i2(intermediate_reg_0[2856]),.o(intermediate_reg_1[1428])); 
fsm fsm_inst_1_372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2855]),.i2(intermediate_reg_0[2854]),.o(intermediate_reg_1[1427])); 
mux_module mux_module_inst_1_373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2853]),.i2(intermediate_reg_0[2852]),.o(intermediate_reg_1[1426]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2851]),.i2(intermediate_reg_0[2850]),.o(intermediate_reg_1[1425]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2849]),.i2(intermediate_reg_0[2848]),.o(intermediate_reg_1[1424])); 
fsm fsm_inst_1_376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2847]),.i2(intermediate_reg_0[2846]),.o(intermediate_reg_1[1423])); 
mux_module mux_module_inst_1_377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2845]),.i2(intermediate_reg_0[2844]),.o(intermediate_reg_1[1422]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2843]),.i2(intermediate_reg_0[2842]),.o(intermediate_reg_1[1421])); 
fsm fsm_inst_1_379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2841]),.i2(intermediate_reg_0[2840]),.o(intermediate_reg_1[1420])); 
fsm fsm_inst_1_380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2839]),.i2(intermediate_reg_0[2838]),.o(intermediate_reg_1[1419])); 
fsm fsm_inst_1_381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2837]),.i2(intermediate_reg_0[2836]),.o(intermediate_reg_1[1418])); 
mux_module mux_module_inst_1_382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2835]),.i2(intermediate_reg_0[2834]),.o(intermediate_reg_1[1417]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2833]),.i2(intermediate_reg_0[2832]),.o(intermediate_reg_1[1416]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2831]),.i2(intermediate_reg_0[2830]),.o(intermediate_reg_1[1415]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2829]),.i2(intermediate_reg_0[2828]),.o(intermediate_reg_1[1414]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2827]),.i2(intermediate_reg_0[2826]),.o(intermediate_reg_1[1413]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2825]),.i2(intermediate_reg_0[2824]),.o(intermediate_reg_1[1412]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2823]),.i2(intermediate_reg_0[2822]),.o(intermediate_reg_1[1411])); 
mux_module mux_module_inst_1_389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2821]),.i2(intermediate_reg_0[2820]),.o(intermediate_reg_1[1410]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2819]),.i2(intermediate_reg_0[2818]),.o(intermediate_reg_1[1409])); 
mux_module mux_module_inst_1_391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2817]),.i2(intermediate_reg_0[2816]),.o(intermediate_reg_1[1408]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2815]),.i2(intermediate_reg_0[2814]),.o(intermediate_reg_1[1407]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2813]),.i2(intermediate_reg_0[2812]),.o(intermediate_reg_1[1406]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2811]),.i2(intermediate_reg_0[2810]),.o(intermediate_reg_1[1405])); 
mux_module mux_module_inst_1_395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2809]),.i2(intermediate_reg_0[2808]),.o(intermediate_reg_1[1404]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2807]),.i2(intermediate_reg_0[2806]),.o(intermediate_reg_1[1403]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2805]),.i2(intermediate_reg_0[2804]),.o(intermediate_reg_1[1402])); 
fsm fsm_inst_1_398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2803]),.i2(intermediate_reg_0[2802]),.o(intermediate_reg_1[1401])); 
fsm fsm_inst_1_399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2801]),.i2(intermediate_reg_0[2800]),.o(intermediate_reg_1[1400])); 
fsm fsm_inst_1_400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2799]),.i2(intermediate_reg_0[2798]),.o(intermediate_reg_1[1399])); 
fsm fsm_inst_1_401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2797]),.i2(intermediate_reg_0[2796]),.o(intermediate_reg_1[1398])); 
fsm fsm_inst_1_402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2795]),.i2(intermediate_reg_0[2794]),.o(intermediate_reg_1[1397])); 
mux_module mux_module_inst_1_403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2793]),.i2(intermediate_reg_0[2792]),.o(intermediate_reg_1[1396]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2791]),.i2(intermediate_reg_0[2790]),.o(intermediate_reg_1[1395]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2789]),.i2(intermediate_reg_0[2788]),.o(intermediate_reg_1[1394])); 
mux_module mux_module_inst_1_406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2787]),.i2(intermediate_reg_0[2786]),.o(intermediate_reg_1[1393]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2785]),.i2(intermediate_reg_0[2784]),.o(intermediate_reg_1[1392]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2783]),.i2(intermediate_reg_0[2782]),.o(intermediate_reg_1[1391])); 
mux_module mux_module_inst_1_409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2781]),.i2(intermediate_reg_0[2780]),.o(intermediate_reg_1[1390]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2779]),.i2(intermediate_reg_0[2778]),.o(intermediate_reg_1[1389]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2777]),.i2(intermediate_reg_0[2776]),.o(intermediate_reg_1[1388]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2775]),.i2(intermediate_reg_0[2774]),.o(intermediate_reg_1[1387]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2773]),.i2(intermediate_reg_0[2772]),.o(intermediate_reg_1[1386]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2771]),.i2(intermediate_reg_0[2770]),.o(intermediate_reg_1[1385]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2769]),.i2(intermediate_reg_0[2768]),.o(intermediate_reg_1[1384])); 
mux_module mux_module_inst_1_416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2767]),.i2(intermediate_reg_0[2766]),.o(intermediate_reg_1[1383]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2765]),.i2(intermediate_reg_0[2764]),.o(intermediate_reg_1[1382])); 
fsm fsm_inst_1_418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2763]),.i2(intermediate_reg_0[2762]),.o(intermediate_reg_1[1381])); 
mux_module mux_module_inst_1_419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2761]),.i2(intermediate_reg_0[2760]),.o(intermediate_reg_1[1380]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2759]),.i2(intermediate_reg_0[2758]),.o(intermediate_reg_1[1379])); 
fsm fsm_inst_1_421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2757]),.i2(intermediate_reg_0[2756]),.o(intermediate_reg_1[1378])); 
mux_module mux_module_inst_1_422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2755]),.i2(intermediate_reg_0[2754]),.o(intermediate_reg_1[1377]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2753]),.i2(intermediate_reg_0[2752]),.o(intermediate_reg_1[1376])); 
fsm fsm_inst_1_424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2751]),.i2(intermediate_reg_0[2750]),.o(intermediate_reg_1[1375])); 
fsm fsm_inst_1_425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2749]),.i2(intermediate_reg_0[2748]),.o(intermediate_reg_1[1374])); 
fsm fsm_inst_1_426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2747]),.i2(intermediate_reg_0[2746]),.o(intermediate_reg_1[1373])); 
mux_module mux_module_inst_1_427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2745]),.i2(intermediate_reg_0[2744]),.o(intermediate_reg_1[1372]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2743]),.i2(intermediate_reg_0[2742]),.o(intermediate_reg_1[1371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2741]),.i2(intermediate_reg_0[2740]),.o(intermediate_reg_1[1370]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2739]),.i2(intermediate_reg_0[2738]),.o(intermediate_reg_1[1369])); 
mux_module mux_module_inst_1_431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2737]),.i2(intermediate_reg_0[2736]),.o(intermediate_reg_1[1368]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2735]),.i2(intermediate_reg_0[2734]),.o(intermediate_reg_1[1367]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2733]),.i2(intermediate_reg_0[2732]),.o(intermediate_reg_1[1366])); 
mux_module mux_module_inst_1_434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2731]),.i2(intermediate_reg_0[2730]),.o(intermediate_reg_1[1365]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2729]),.i2(intermediate_reg_0[2728]),.o(intermediate_reg_1[1364])); 
mux_module mux_module_inst_1_436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2727]),.i2(intermediate_reg_0[2726]),.o(intermediate_reg_1[1363]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2725]),.i2(intermediate_reg_0[2724]),.o(intermediate_reg_1[1362])); 
mux_module mux_module_inst_1_438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2723]),.i2(intermediate_reg_0[2722]),.o(intermediate_reg_1[1361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2721]),.i2(intermediate_reg_0[2720]),.o(intermediate_reg_1[1360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2719]),.i2(intermediate_reg_0[2718]),.o(intermediate_reg_1[1359]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2717]),.i2(intermediate_reg_0[2716]),.o(intermediate_reg_1[1358])); 
mux_module mux_module_inst_1_442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2715]),.i2(intermediate_reg_0[2714]),.o(intermediate_reg_1[1357]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2713]),.i2(intermediate_reg_0[2712]),.o(intermediate_reg_1[1356]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2711]),.i2(intermediate_reg_0[2710]),.o(intermediate_reg_1[1355]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2709]),.i2(intermediate_reg_0[2708]),.o(intermediate_reg_1[1354])); 
mux_module mux_module_inst_1_446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2707]),.i2(intermediate_reg_0[2706]),.o(intermediate_reg_1[1353]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2705]),.i2(intermediate_reg_0[2704]),.o(intermediate_reg_1[1352])); 
mux_module mux_module_inst_1_448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2703]),.i2(intermediate_reg_0[2702]),.o(intermediate_reg_1[1351]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2701]),.i2(intermediate_reg_0[2700]),.o(intermediate_reg_1[1350])); 
fsm fsm_inst_1_450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2699]),.i2(intermediate_reg_0[2698]),.o(intermediate_reg_1[1349])); 
fsm fsm_inst_1_451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2697]),.i2(intermediate_reg_0[2696]),.o(intermediate_reg_1[1348])); 
mux_module mux_module_inst_1_452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2695]),.i2(intermediate_reg_0[2694]),.o(intermediate_reg_1[1347]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2693]),.i2(intermediate_reg_0[2692]),.o(intermediate_reg_1[1346])); 
fsm fsm_inst_1_454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2691]),.i2(intermediate_reg_0[2690]),.o(intermediate_reg_1[1345])); 
fsm fsm_inst_1_455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2689]),.i2(intermediate_reg_0[2688]),.o(intermediate_reg_1[1344])); 
fsm fsm_inst_1_456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2687]),.i2(intermediate_reg_0[2686]),.o(intermediate_reg_1[1343])); 
fsm fsm_inst_1_457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2685]),.i2(intermediate_reg_0[2684]),.o(intermediate_reg_1[1342])); 
fsm fsm_inst_1_458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2683]),.i2(intermediate_reg_0[2682]),.o(intermediate_reg_1[1341])); 
mux_module mux_module_inst_1_459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2681]),.i2(intermediate_reg_0[2680]),.o(intermediate_reg_1[1340]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2679]),.i2(intermediate_reg_0[2678]),.o(intermediate_reg_1[1339]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2677]),.i2(intermediate_reg_0[2676]),.o(intermediate_reg_1[1338])); 
fsm fsm_inst_1_462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2675]),.i2(intermediate_reg_0[2674]),.o(intermediate_reg_1[1337])); 
mux_module mux_module_inst_1_463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2673]),.i2(intermediate_reg_0[2672]),.o(intermediate_reg_1[1336]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2671]),.i2(intermediate_reg_0[2670]),.o(intermediate_reg_1[1335]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2669]),.i2(intermediate_reg_0[2668]),.o(intermediate_reg_1[1334]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2667]),.i2(intermediate_reg_0[2666]),.o(intermediate_reg_1[1333])); 
mux_module mux_module_inst_1_467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2665]),.i2(intermediate_reg_0[2664]),.o(intermediate_reg_1[1332]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2663]),.i2(intermediate_reg_0[2662]),.o(intermediate_reg_1[1331])); 
mux_module mux_module_inst_1_469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2661]),.i2(intermediate_reg_0[2660]),.o(intermediate_reg_1[1330]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2659]),.i2(intermediate_reg_0[2658]),.o(intermediate_reg_1[1329])); 
mux_module mux_module_inst_1_471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2657]),.i2(intermediate_reg_0[2656]),.o(intermediate_reg_1[1328]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2655]),.i2(intermediate_reg_0[2654]),.o(intermediate_reg_1[1327])); 
fsm fsm_inst_1_473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2653]),.i2(intermediate_reg_0[2652]),.o(intermediate_reg_1[1326])); 
fsm fsm_inst_1_474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2651]),.i2(intermediate_reg_0[2650]),.o(intermediate_reg_1[1325])); 
fsm fsm_inst_1_475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2649]),.i2(intermediate_reg_0[2648]),.o(intermediate_reg_1[1324])); 
fsm fsm_inst_1_476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2647]),.i2(intermediate_reg_0[2646]),.o(intermediate_reg_1[1323])); 
fsm fsm_inst_1_477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2645]),.i2(intermediate_reg_0[2644]),.o(intermediate_reg_1[1322])); 
mux_module mux_module_inst_1_478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2643]),.i2(intermediate_reg_0[2642]),.o(intermediate_reg_1[1321]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2641]),.i2(intermediate_reg_0[2640]),.o(intermediate_reg_1[1320])); 
fsm fsm_inst_1_480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2639]),.i2(intermediate_reg_0[2638]),.o(intermediate_reg_1[1319])); 
fsm fsm_inst_1_481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2637]),.i2(intermediate_reg_0[2636]),.o(intermediate_reg_1[1318])); 
mux_module mux_module_inst_1_482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2635]),.i2(intermediate_reg_0[2634]),.o(intermediate_reg_1[1317]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2633]),.i2(intermediate_reg_0[2632]),.o(intermediate_reg_1[1316])); 
mux_module mux_module_inst_1_484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2631]),.i2(intermediate_reg_0[2630]),.o(intermediate_reg_1[1315]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2629]),.i2(intermediate_reg_0[2628]),.o(intermediate_reg_1[1314])); 
mux_module mux_module_inst_1_486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2627]),.i2(intermediate_reg_0[2626]),.o(intermediate_reg_1[1313]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2625]),.i2(intermediate_reg_0[2624]),.o(intermediate_reg_1[1312]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2623]),.i2(intermediate_reg_0[2622]),.o(intermediate_reg_1[1311])); 
fsm fsm_inst_1_489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2621]),.i2(intermediate_reg_0[2620]),.o(intermediate_reg_1[1310])); 
mux_module mux_module_inst_1_490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2619]),.i2(intermediate_reg_0[2618]),.o(intermediate_reg_1[1309]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2617]),.i2(intermediate_reg_0[2616]),.o(intermediate_reg_1[1308])); 
fsm fsm_inst_1_492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2615]),.i2(intermediate_reg_0[2614]),.o(intermediate_reg_1[1307])); 
fsm fsm_inst_1_493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2613]),.i2(intermediate_reg_0[2612]),.o(intermediate_reg_1[1306])); 
mux_module mux_module_inst_1_494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2611]),.i2(intermediate_reg_0[2610]),.o(intermediate_reg_1[1305]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2609]),.i2(intermediate_reg_0[2608]),.o(intermediate_reg_1[1304])); 
mux_module mux_module_inst_1_496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2607]),.i2(intermediate_reg_0[2606]),.o(intermediate_reg_1[1303]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2605]),.i2(intermediate_reg_0[2604]),.o(intermediate_reg_1[1302]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2603]),.i2(intermediate_reg_0[2602]),.o(intermediate_reg_1[1301]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2601]),.i2(intermediate_reg_0[2600]),.o(intermediate_reg_1[1300])); 
fsm fsm_inst_1_500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2599]),.i2(intermediate_reg_0[2598]),.o(intermediate_reg_1[1299])); 
mux_module mux_module_inst_1_501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2597]),.i2(intermediate_reg_0[2596]),.o(intermediate_reg_1[1298]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2595]),.i2(intermediate_reg_0[2594]),.o(intermediate_reg_1[1297]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2593]),.i2(intermediate_reg_0[2592]),.o(intermediate_reg_1[1296])); 
fsm fsm_inst_1_504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2591]),.i2(intermediate_reg_0[2590]),.o(intermediate_reg_1[1295])); 
fsm fsm_inst_1_505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2589]),.i2(intermediate_reg_0[2588]),.o(intermediate_reg_1[1294])); 
fsm fsm_inst_1_506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2587]),.i2(intermediate_reg_0[2586]),.o(intermediate_reg_1[1293])); 
mux_module mux_module_inst_1_507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2585]),.i2(intermediate_reg_0[2584]),.o(intermediate_reg_1[1292]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2583]),.i2(intermediate_reg_0[2582]),.o(intermediate_reg_1[1291]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2581]),.i2(intermediate_reg_0[2580]),.o(intermediate_reg_1[1290]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2579]),.i2(intermediate_reg_0[2578]),.o(intermediate_reg_1[1289])); 
fsm fsm_inst_1_511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2577]),.i2(intermediate_reg_0[2576]),.o(intermediate_reg_1[1288])); 
fsm fsm_inst_1_512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2575]),.i2(intermediate_reg_0[2574]),.o(intermediate_reg_1[1287])); 
fsm fsm_inst_1_513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2573]),.i2(intermediate_reg_0[2572]),.o(intermediate_reg_1[1286])); 
mux_module mux_module_inst_1_514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2571]),.i2(intermediate_reg_0[2570]),.o(intermediate_reg_1[1285]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2569]),.i2(intermediate_reg_0[2568]),.o(intermediate_reg_1[1284])); 
mux_module mux_module_inst_1_516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2567]),.i2(intermediate_reg_0[2566]),.o(intermediate_reg_1[1283]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2565]),.i2(intermediate_reg_0[2564]),.o(intermediate_reg_1[1282])); 
fsm fsm_inst_1_518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2563]),.i2(intermediate_reg_0[2562]),.o(intermediate_reg_1[1281])); 
fsm fsm_inst_1_519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2561]),.i2(intermediate_reg_0[2560]),.o(intermediate_reg_1[1280])); 
mux_module mux_module_inst_1_520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2559]),.i2(intermediate_reg_0[2558]),.o(intermediate_reg_1[1279]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2557]),.i2(intermediate_reg_0[2556]),.o(intermediate_reg_1[1278])); 
mux_module mux_module_inst_1_522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2555]),.i2(intermediate_reg_0[2554]),.o(intermediate_reg_1[1277]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2553]),.i2(intermediate_reg_0[2552]),.o(intermediate_reg_1[1276]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2551]),.i2(intermediate_reg_0[2550]),.o(intermediate_reg_1[1275]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2549]),.i2(intermediate_reg_0[2548]),.o(intermediate_reg_1[1274]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2547]),.i2(intermediate_reg_0[2546]),.o(intermediate_reg_1[1273])); 
fsm fsm_inst_1_527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2545]),.i2(intermediate_reg_0[2544]),.o(intermediate_reg_1[1272])); 
fsm fsm_inst_1_528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2543]),.i2(intermediate_reg_0[2542]),.o(intermediate_reg_1[1271])); 
mux_module mux_module_inst_1_529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2541]),.i2(intermediate_reg_0[2540]),.o(intermediate_reg_1[1270]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2539]),.i2(intermediate_reg_0[2538]),.o(intermediate_reg_1[1269]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2537]),.i2(intermediate_reg_0[2536]),.o(intermediate_reg_1[1268])); 
mux_module mux_module_inst_1_532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2535]),.i2(intermediate_reg_0[2534]),.o(intermediate_reg_1[1267]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2533]),.i2(intermediate_reg_0[2532]),.o(intermediate_reg_1[1266])); 
mux_module mux_module_inst_1_534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2531]),.i2(intermediate_reg_0[2530]),.o(intermediate_reg_1[1265]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2529]),.i2(intermediate_reg_0[2528]),.o(intermediate_reg_1[1264]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2527]),.i2(intermediate_reg_0[2526]),.o(intermediate_reg_1[1263]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2525]),.i2(intermediate_reg_0[2524]),.o(intermediate_reg_1[1262]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2523]),.i2(intermediate_reg_0[2522]),.o(intermediate_reg_1[1261]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2521]),.i2(intermediate_reg_0[2520]),.o(intermediate_reg_1[1260]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2519]),.i2(intermediate_reg_0[2518]),.o(intermediate_reg_1[1259])); 
fsm fsm_inst_1_541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2517]),.i2(intermediate_reg_0[2516]),.o(intermediate_reg_1[1258])); 
fsm fsm_inst_1_542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2515]),.i2(intermediate_reg_0[2514]),.o(intermediate_reg_1[1257])); 
fsm fsm_inst_1_543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2513]),.i2(intermediate_reg_0[2512]),.o(intermediate_reg_1[1256])); 
fsm fsm_inst_1_544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2511]),.i2(intermediate_reg_0[2510]),.o(intermediate_reg_1[1255])); 
fsm fsm_inst_1_545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2509]),.i2(intermediate_reg_0[2508]),.o(intermediate_reg_1[1254])); 
fsm fsm_inst_1_546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2507]),.i2(intermediate_reg_0[2506]),.o(intermediate_reg_1[1253])); 
mux_module mux_module_inst_1_547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2505]),.i2(intermediate_reg_0[2504]),.o(intermediate_reg_1[1252]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2503]),.i2(intermediate_reg_0[2502]),.o(intermediate_reg_1[1251]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2501]),.i2(intermediate_reg_0[2500]),.o(intermediate_reg_1[1250])); 
fsm fsm_inst_1_550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2499]),.i2(intermediate_reg_0[2498]),.o(intermediate_reg_1[1249])); 
mux_module mux_module_inst_1_551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2497]),.i2(intermediate_reg_0[2496]),.o(intermediate_reg_1[1248]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2495]),.i2(intermediate_reg_0[2494]),.o(intermediate_reg_1[1247]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2493]),.i2(intermediate_reg_0[2492]),.o(intermediate_reg_1[1246])); 
fsm fsm_inst_1_554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2491]),.i2(intermediate_reg_0[2490]),.o(intermediate_reg_1[1245])); 
mux_module mux_module_inst_1_555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2489]),.i2(intermediate_reg_0[2488]),.o(intermediate_reg_1[1244]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2487]),.i2(intermediate_reg_0[2486]),.o(intermediate_reg_1[1243])); 
mux_module mux_module_inst_1_557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2485]),.i2(intermediate_reg_0[2484]),.o(intermediate_reg_1[1242]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2483]),.i2(intermediate_reg_0[2482]),.o(intermediate_reg_1[1241]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2481]),.i2(intermediate_reg_0[2480]),.o(intermediate_reg_1[1240])); 
mux_module mux_module_inst_1_560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2479]),.i2(intermediate_reg_0[2478]),.o(intermediate_reg_1[1239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2477]),.i2(intermediate_reg_0[2476]),.o(intermediate_reg_1[1238]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2475]),.i2(intermediate_reg_0[2474]),.o(intermediate_reg_1[1237])); 
fsm fsm_inst_1_563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2473]),.i2(intermediate_reg_0[2472]),.o(intermediate_reg_1[1236])); 
mux_module mux_module_inst_1_564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2471]),.i2(intermediate_reg_0[2470]),.o(intermediate_reg_1[1235]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2469]),.i2(intermediate_reg_0[2468]),.o(intermediate_reg_1[1234]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2467]),.i2(intermediate_reg_0[2466]),.o(intermediate_reg_1[1233]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2465]),.i2(intermediate_reg_0[2464]),.o(intermediate_reg_1[1232])); 
fsm fsm_inst_1_568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2463]),.i2(intermediate_reg_0[2462]),.o(intermediate_reg_1[1231])); 
mux_module mux_module_inst_1_569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2461]),.i2(intermediate_reg_0[2460]),.o(intermediate_reg_1[1230]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2459]),.i2(intermediate_reg_0[2458]),.o(intermediate_reg_1[1229]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2457]),.i2(intermediate_reg_0[2456]),.o(intermediate_reg_1[1228]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2455]),.i2(intermediate_reg_0[2454]),.o(intermediate_reg_1[1227]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2453]),.i2(intermediate_reg_0[2452]),.o(intermediate_reg_1[1226])); 
fsm fsm_inst_1_574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2451]),.i2(intermediate_reg_0[2450]),.o(intermediate_reg_1[1225])); 
mux_module mux_module_inst_1_575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2449]),.i2(intermediate_reg_0[2448]),.o(intermediate_reg_1[1224]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2447]),.i2(intermediate_reg_0[2446]),.o(intermediate_reg_1[1223]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2445]),.i2(intermediate_reg_0[2444]),.o(intermediate_reg_1[1222]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2443]),.i2(intermediate_reg_0[2442]),.o(intermediate_reg_1[1221]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2441]),.i2(intermediate_reg_0[2440]),.o(intermediate_reg_1[1220])); 
fsm fsm_inst_1_580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2439]),.i2(intermediate_reg_0[2438]),.o(intermediate_reg_1[1219])); 
mux_module mux_module_inst_1_581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2437]),.i2(intermediate_reg_0[2436]),.o(intermediate_reg_1[1218]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2435]),.i2(intermediate_reg_0[2434]),.o(intermediate_reg_1[1217])); 
fsm fsm_inst_1_583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2433]),.i2(intermediate_reg_0[2432]),.o(intermediate_reg_1[1216])); 
fsm fsm_inst_1_584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2431]),.i2(intermediate_reg_0[2430]),.o(intermediate_reg_1[1215])); 
fsm fsm_inst_1_585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2429]),.i2(intermediate_reg_0[2428]),.o(intermediate_reg_1[1214])); 
mux_module mux_module_inst_1_586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2427]),.i2(intermediate_reg_0[2426]),.o(intermediate_reg_1[1213]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2425]),.i2(intermediate_reg_0[2424]),.o(intermediate_reg_1[1212])); 
mux_module mux_module_inst_1_588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2423]),.i2(intermediate_reg_0[2422]),.o(intermediate_reg_1[1211]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2421]),.i2(intermediate_reg_0[2420]),.o(intermediate_reg_1[1210])); 
fsm fsm_inst_1_590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2419]),.i2(intermediate_reg_0[2418]),.o(intermediate_reg_1[1209])); 
fsm fsm_inst_1_591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2417]),.i2(intermediate_reg_0[2416]),.o(intermediate_reg_1[1208])); 
fsm fsm_inst_1_592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2415]),.i2(intermediate_reg_0[2414]),.o(intermediate_reg_1[1207])); 
fsm fsm_inst_1_593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2413]),.i2(intermediate_reg_0[2412]),.o(intermediate_reg_1[1206])); 
fsm fsm_inst_1_594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2411]),.i2(intermediate_reg_0[2410]),.o(intermediate_reg_1[1205])); 
mux_module mux_module_inst_1_595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2409]),.i2(intermediate_reg_0[2408]),.o(intermediate_reg_1[1204]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2407]),.i2(intermediate_reg_0[2406]),.o(intermediate_reg_1[1203]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2405]),.i2(intermediate_reg_0[2404]),.o(intermediate_reg_1[1202])); 
fsm fsm_inst_1_598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2403]),.i2(intermediate_reg_0[2402]),.o(intermediate_reg_1[1201])); 
mux_module mux_module_inst_1_599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2401]),.i2(intermediate_reg_0[2400]),.o(intermediate_reg_1[1200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2399]),.i2(intermediate_reg_0[2398]),.o(intermediate_reg_1[1199]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2397]),.i2(intermediate_reg_0[2396]),.o(intermediate_reg_1[1198])); 
fsm fsm_inst_1_602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2395]),.i2(intermediate_reg_0[2394]),.o(intermediate_reg_1[1197])); 
mux_module mux_module_inst_1_603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2393]),.i2(intermediate_reg_0[2392]),.o(intermediate_reg_1[1196]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2391]),.i2(intermediate_reg_0[2390]),.o(intermediate_reg_1[1195])); 
mux_module mux_module_inst_1_605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2389]),.i2(intermediate_reg_0[2388]),.o(intermediate_reg_1[1194]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2387]),.i2(intermediate_reg_0[2386]),.o(intermediate_reg_1[1193])); 
mux_module mux_module_inst_1_607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2385]),.i2(intermediate_reg_0[2384]),.o(intermediate_reg_1[1192]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2383]),.i2(intermediate_reg_0[2382]),.o(intermediate_reg_1[1191]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2381]),.i2(intermediate_reg_0[2380]),.o(intermediate_reg_1[1190])); 
mux_module mux_module_inst_1_610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2379]),.i2(intermediate_reg_0[2378]),.o(intermediate_reg_1[1189]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2377]),.i2(intermediate_reg_0[2376]),.o(intermediate_reg_1[1188]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2375]),.i2(intermediate_reg_0[2374]),.o(intermediate_reg_1[1187]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2373]),.i2(intermediate_reg_0[2372]),.o(intermediate_reg_1[1186])); 
mux_module mux_module_inst_1_614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2371]),.i2(intermediate_reg_0[2370]),.o(intermediate_reg_1[1185]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2369]),.i2(intermediate_reg_0[2368]),.o(intermediate_reg_1[1184]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2367]),.i2(intermediate_reg_0[2366]),.o(intermediate_reg_1[1183])); 
mux_module mux_module_inst_1_617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2365]),.i2(intermediate_reg_0[2364]),.o(intermediate_reg_1[1182]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2363]),.i2(intermediate_reg_0[2362]),.o(intermediate_reg_1[1181])); 
fsm fsm_inst_1_619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2361]),.i2(intermediate_reg_0[2360]),.o(intermediate_reg_1[1180])); 
mux_module mux_module_inst_1_620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2359]),.i2(intermediate_reg_0[2358]),.o(intermediate_reg_1[1179]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2357]),.i2(intermediate_reg_0[2356]),.o(intermediate_reg_1[1178]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2355]),.i2(intermediate_reg_0[2354]),.o(intermediate_reg_1[1177]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2353]),.i2(intermediate_reg_0[2352]),.o(intermediate_reg_1[1176])); 
fsm fsm_inst_1_624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2351]),.i2(intermediate_reg_0[2350]),.o(intermediate_reg_1[1175])); 
fsm fsm_inst_1_625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2349]),.i2(intermediate_reg_0[2348]),.o(intermediate_reg_1[1174])); 
mux_module mux_module_inst_1_626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2347]),.i2(intermediate_reg_0[2346]),.o(intermediate_reg_1[1173]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2345]),.i2(intermediate_reg_0[2344]),.o(intermediate_reg_1[1172]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2343]),.i2(intermediate_reg_0[2342]),.o(intermediate_reg_1[1171])); 
mux_module mux_module_inst_1_629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2341]),.i2(intermediate_reg_0[2340]),.o(intermediate_reg_1[1170]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2339]),.i2(intermediate_reg_0[2338]),.o(intermediate_reg_1[1169])); 
fsm fsm_inst_1_631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2337]),.i2(intermediate_reg_0[2336]),.o(intermediate_reg_1[1168])); 
mux_module mux_module_inst_1_632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2335]),.i2(intermediate_reg_0[2334]),.o(intermediate_reg_1[1167]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2333]),.i2(intermediate_reg_0[2332]),.o(intermediate_reg_1[1166]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2331]),.i2(intermediate_reg_0[2330]),.o(intermediate_reg_1[1165])); 
fsm fsm_inst_1_635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2329]),.i2(intermediate_reg_0[2328]),.o(intermediate_reg_1[1164])); 
fsm fsm_inst_1_636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2327]),.i2(intermediate_reg_0[2326]),.o(intermediate_reg_1[1163])); 
fsm fsm_inst_1_637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2325]),.i2(intermediate_reg_0[2324]),.o(intermediate_reg_1[1162])); 
mux_module mux_module_inst_1_638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2323]),.i2(intermediate_reg_0[2322]),.o(intermediate_reg_1[1161]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2321]),.i2(intermediate_reg_0[2320]),.o(intermediate_reg_1[1160])); 
mux_module mux_module_inst_1_640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2319]),.i2(intermediate_reg_0[2318]),.o(intermediate_reg_1[1159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2317]),.i2(intermediate_reg_0[2316]),.o(intermediate_reg_1[1158]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2315]),.i2(intermediate_reg_0[2314]),.o(intermediate_reg_1[1157])); 
fsm fsm_inst_1_643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2313]),.i2(intermediate_reg_0[2312]),.o(intermediate_reg_1[1156])); 
fsm fsm_inst_1_644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2311]),.i2(intermediate_reg_0[2310]),.o(intermediate_reg_1[1155])); 
mux_module mux_module_inst_1_645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2309]),.i2(intermediate_reg_0[2308]),.o(intermediate_reg_1[1154]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2307]),.i2(intermediate_reg_0[2306]),.o(intermediate_reg_1[1153]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2305]),.i2(intermediate_reg_0[2304]),.o(intermediate_reg_1[1152]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2303]),.i2(intermediate_reg_0[2302]),.o(intermediate_reg_1[1151]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2301]),.i2(intermediate_reg_0[2300]),.o(intermediate_reg_1[1150]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2299]),.i2(intermediate_reg_0[2298]),.o(intermediate_reg_1[1149])); 
fsm fsm_inst_1_651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2297]),.i2(intermediate_reg_0[2296]),.o(intermediate_reg_1[1148])); 
fsm fsm_inst_1_652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2295]),.i2(intermediate_reg_0[2294]),.o(intermediate_reg_1[1147])); 
mux_module mux_module_inst_1_653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2293]),.i2(intermediate_reg_0[2292]),.o(intermediate_reg_1[1146]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2291]),.i2(intermediate_reg_0[2290]),.o(intermediate_reg_1[1145]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2289]),.i2(intermediate_reg_0[2288]),.o(intermediate_reg_1[1144]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2287]),.i2(intermediate_reg_0[2286]),.o(intermediate_reg_1[1143]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2285]),.i2(intermediate_reg_0[2284]),.o(intermediate_reg_1[1142]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2283]),.i2(intermediate_reg_0[2282]),.o(intermediate_reg_1[1141]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2281]),.i2(intermediate_reg_0[2280]),.o(intermediate_reg_1[1140])); 
mux_module mux_module_inst_1_660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2279]),.i2(intermediate_reg_0[2278]),.o(intermediate_reg_1[1139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2277]),.i2(intermediate_reg_0[2276]),.o(intermediate_reg_1[1138]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2275]),.i2(intermediate_reg_0[2274]),.o(intermediate_reg_1[1137])); 
fsm fsm_inst_1_663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2273]),.i2(intermediate_reg_0[2272]),.o(intermediate_reg_1[1136])); 
mux_module mux_module_inst_1_664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2271]),.i2(intermediate_reg_0[2270]),.o(intermediate_reg_1[1135]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2269]),.i2(intermediate_reg_0[2268]),.o(intermediate_reg_1[1134])); 
mux_module mux_module_inst_1_666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2267]),.i2(intermediate_reg_0[2266]),.o(intermediate_reg_1[1133]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2265]),.i2(intermediate_reg_0[2264]),.o(intermediate_reg_1[1132])); 
mux_module mux_module_inst_1_668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2263]),.i2(intermediate_reg_0[2262]),.o(intermediate_reg_1[1131]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2261]),.i2(intermediate_reg_0[2260]),.o(intermediate_reg_1[1130])); 
fsm fsm_inst_1_670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2259]),.i2(intermediate_reg_0[2258]),.o(intermediate_reg_1[1129])); 
mux_module mux_module_inst_1_671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2257]),.i2(intermediate_reg_0[2256]),.o(intermediate_reg_1[1128]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2255]),.i2(intermediate_reg_0[2254]),.o(intermediate_reg_1[1127]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2253]),.i2(intermediate_reg_0[2252]),.o(intermediate_reg_1[1126])); 
fsm fsm_inst_1_674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2251]),.i2(intermediate_reg_0[2250]),.o(intermediate_reg_1[1125])); 
fsm fsm_inst_1_675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2249]),.i2(intermediate_reg_0[2248]),.o(intermediate_reg_1[1124])); 
fsm fsm_inst_1_676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2247]),.i2(intermediate_reg_0[2246]),.o(intermediate_reg_1[1123])); 
fsm fsm_inst_1_677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2245]),.i2(intermediate_reg_0[2244]),.o(intermediate_reg_1[1122])); 
fsm fsm_inst_1_678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2243]),.i2(intermediate_reg_0[2242]),.o(intermediate_reg_1[1121])); 
fsm fsm_inst_1_679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2241]),.i2(intermediate_reg_0[2240]),.o(intermediate_reg_1[1120])); 
mux_module mux_module_inst_1_680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2239]),.i2(intermediate_reg_0[2238]),.o(intermediate_reg_1[1119]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2237]),.i2(intermediate_reg_0[2236]),.o(intermediate_reg_1[1118])); 
mux_module mux_module_inst_1_682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2235]),.i2(intermediate_reg_0[2234]),.o(intermediate_reg_1[1117]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2233]),.i2(intermediate_reg_0[2232]),.o(intermediate_reg_1[1116])); 
mux_module mux_module_inst_1_684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2231]),.i2(intermediate_reg_0[2230]),.o(intermediate_reg_1[1115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2229]),.i2(intermediate_reg_0[2228]),.o(intermediate_reg_1[1114])); 
mux_module mux_module_inst_1_686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2227]),.i2(intermediate_reg_0[2226]),.o(intermediate_reg_1[1113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2225]),.i2(intermediate_reg_0[2224]),.o(intermediate_reg_1[1112]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2223]),.i2(intermediate_reg_0[2222]),.o(intermediate_reg_1[1111])); 
mux_module mux_module_inst_1_689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2221]),.i2(intermediate_reg_0[2220]),.o(intermediate_reg_1[1110]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2219]),.i2(intermediate_reg_0[2218]),.o(intermediate_reg_1[1109]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2217]),.i2(intermediate_reg_0[2216]),.o(intermediate_reg_1[1108])); 
fsm fsm_inst_1_692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2215]),.i2(intermediate_reg_0[2214]),.o(intermediate_reg_1[1107])); 
mux_module mux_module_inst_1_693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2213]),.i2(intermediate_reg_0[2212]),.o(intermediate_reg_1[1106]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2211]),.i2(intermediate_reg_0[2210]),.o(intermediate_reg_1[1105])); 
fsm fsm_inst_1_695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2209]),.i2(intermediate_reg_0[2208]),.o(intermediate_reg_1[1104])); 
fsm fsm_inst_1_696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2207]),.i2(intermediate_reg_0[2206]),.o(intermediate_reg_1[1103])); 
mux_module mux_module_inst_1_697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2205]),.i2(intermediate_reg_0[2204]),.o(intermediate_reg_1[1102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2203]),.i2(intermediate_reg_0[2202]),.o(intermediate_reg_1[1101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2201]),.i2(intermediate_reg_0[2200]),.o(intermediate_reg_1[1100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2199]),.i2(intermediate_reg_0[2198]),.o(intermediate_reg_1[1099]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2197]),.i2(intermediate_reg_0[2196]),.o(intermediate_reg_1[1098]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2195]),.i2(intermediate_reg_0[2194]),.o(intermediate_reg_1[1097]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2193]),.i2(intermediate_reg_0[2192]),.o(intermediate_reg_1[1096])); 
mux_module mux_module_inst_1_704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2191]),.i2(intermediate_reg_0[2190]),.o(intermediate_reg_1[1095]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2189]),.i2(intermediate_reg_0[2188]),.o(intermediate_reg_1[1094]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2187]),.i2(intermediate_reg_0[2186]),.o(intermediate_reg_1[1093])); 
mux_module mux_module_inst_1_707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2185]),.i2(intermediate_reg_0[2184]),.o(intermediate_reg_1[1092]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2183]),.i2(intermediate_reg_0[2182]),.o(intermediate_reg_1[1091])); 
fsm fsm_inst_1_709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2181]),.i2(intermediate_reg_0[2180]),.o(intermediate_reg_1[1090])); 
fsm fsm_inst_1_710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2179]),.i2(intermediate_reg_0[2178]),.o(intermediate_reg_1[1089])); 
mux_module mux_module_inst_1_711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2177]),.i2(intermediate_reg_0[2176]),.o(intermediate_reg_1[1088]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2175]),.i2(intermediate_reg_0[2174]),.o(intermediate_reg_1[1087]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2173]),.i2(intermediate_reg_0[2172]),.o(intermediate_reg_1[1086]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2171]),.i2(intermediate_reg_0[2170]),.o(intermediate_reg_1[1085]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2169]),.i2(intermediate_reg_0[2168]),.o(intermediate_reg_1[1084]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2167]),.i2(intermediate_reg_0[2166]),.o(intermediate_reg_1[1083])); 
fsm fsm_inst_1_717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2165]),.i2(intermediate_reg_0[2164]),.o(intermediate_reg_1[1082])); 
mux_module mux_module_inst_1_718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2163]),.i2(intermediate_reg_0[2162]),.o(intermediate_reg_1[1081]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2161]),.i2(intermediate_reg_0[2160]),.o(intermediate_reg_1[1080])); 
mux_module mux_module_inst_1_720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2159]),.i2(intermediate_reg_0[2158]),.o(intermediate_reg_1[1079]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2157]),.i2(intermediate_reg_0[2156]),.o(intermediate_reg_1[1078]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2155]),.i2(intermediate_reg_0[2154]),.o(intermediate_reg_1[1077])); 
mux_module mux_module_inst_1_723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2153]),.i2(intermediate_reg_0[2152]),.o(intermediate_reg_1[1076]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2151]),.i2(intermediate_reg_0[2150]),.o(intermediate_reg_1[1075]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2149]),.i2(intermediate_reg_0[2148]),.o(intermediate_reg_1[1074])); 
fsm fsm_inst_1_726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2147]),.i2(intermediate_reg_0[2146]),.o(intermediate_reg_1[1073])); 
mux_module mux_module_inst_1_727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2145]),.i2(intermediate_reg_0[2144]),.o(intermediate_reg_1[1072]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2143]),.i2(intermediate_reg_0[2142]),.o(intermediate_reg_1[1071]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2141]),.i2(intermediate_reg_0[2140]),.o(intermediate_reg_1[1070])); 
mux_module mux_module_inst_1_730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2139]),.i2(intermediate_reg_0[2138]),.o(intermediate_reg_1[1069]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2137]),.i2(intermediate_reg_0[2136]),.o(intermediate_reg_1[1068]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2135]),.i2(intermediate_reg_0[2134]),.o(intermediate_reg_1[1067])); 
mux_module mux_module_inst_1_733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2133]),.i2(intermediate_reg_0[2132]),.o(intermediate_reg_1[1066]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2131]),.i2(intermediate_reg_0[2130]),.o(intermediate_reg_1[1065])); 
mux_module mux_module_inst_1_735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2129]),.i2(intermediate_reg_0[2128]),.o(intermediate_reg_1[1064]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2127]),.i2(intermediate_reg_0[2126]),.o(intermediate_reg_1[1063]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2125]),.i2(intermediate_reg_0[2124]),.o(intermediate_reg_1[1062]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2123]),.i2(intermediate_reg_0[2122]),.o(intermediate_reg_1[1061]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2121]),.i2(intermediate_reg_0[2120]),.o(intermediate_reg_1[1060]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2119]),.i2(intermediate_reg_0[2118]),.o(intermediate_reg_1[1059])); 
fsm fsm_inst_1_741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2117]),.i2(intermediate_reg_0[2116]),.o(intermediate_reg_1[1058])); 
mux_module mux_module_inst_1_742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2115]),.i2(intermediate_reg_0[2114]),.o(intermediate_reg_1[1057]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2113]),.i2(intermediate_reg_0[2112]),.o(intermediate_reg_1[1056]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2111]),.i2(intermediate_reg_0[2110]),.o(intermediate_reg_1[1055]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2109]),.i2(intermediate_reg_0[2108]),.o(intermediate_reg_1[1054]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2107]),.i2(intermediate_reg_0[2106]),.o(intermediate_reg_1[1053])); 
mux_module mux_module_inst_1_747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2105]),.i2(intermediate_reg_0[2104]),.o(intermediate_reg_1[1052]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2103]),.i2(intermediate_reg_0[2102]),.o(intermediate_reg_1[1051]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2101]),.i2(intermediate_reg_0[2100]),.o(intermediate_reg_1[1050]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2099]),.i2(intermediate_reg_0[2098]),.o(intermediate_reg_1[1049])); 
fsm fsm_inst_1_751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2097]),.i2(intermediate_reg_0[2096]),.o(intermediate_reg_1[1048])); 
mux_module mux_module_inst_1_752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2095]),.i2(intermediate_reg_0[2094]),.o(intermediate_reg_1[1047]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2093]),.i2(intermediate_reg_0[2092]),.o(intermediate_reg_1[1046]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2091]),.i2(intermediate_reg_0[2090]),.o(intermediate_reg_1[1045]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2089]),.i2(intermediate_reg_0[2088]),.o(intermediate_reg_1[1044]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2087]),.i2(intermediate_reg_0[2086]),.o(intermediate_reg_1[1043])); 
fsm fsm_inst_1_757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2085]),.i2(intermediate_reg_0[2084]),.o(intermediate_reg_1[1042])); 
mux_module mux_module_inst_1_758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2083]),.i2(intermediate_reg_0[2082]),.o(intermediate_reg_1[1041]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2081]),.i2(intermediate_reg_0[2080]),.o(intermediate_reg_1[1040])); 
fsm fsm_inst_1_760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2079]),.i2(intermediate_reg_0[2078]),.o(intermediate_reg_1[1039])); 
fsm fsm_inst_1_761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2077]),.i2(intermediate_reg_0[2076]),.o(intermediate_reg_1[1038])); 
fsm fsm_inst_1_762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2075]),.i2(intermediate_reg_0[2074]),.o(intermediate_reg_1[1037])); 
mux_module mux_module_inst_1_763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2073]),.i2(intermediate_reg_0[2072]),.o(intermediate_reg_1[1036]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2071]),.i2(intermediate_reg_0[2070]),.o(intermediate_reg_1[1035]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2069]),.i2(intermediate_reg_0[2068]),.o(intermediate_reg_1[1034]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2067]),.i2(intermediate_reg_0[2066]),.o(intermediate_reg_1[1033]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2065]),.i2(intermediate_reg_0[2064]),.o(intermediate_reg_1[1032]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2063]),.i2(intermediate_reg_0[2062]),.o(intermediate_reg_1[1031]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2061]),.i2(intermediate_reg_0[2060]),.o(intermediate_reg_1[1030])); 
mux_module mux_module_inst_1_770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2059]),.i2(intermediate_reg_0[2058]),.o(intermediate_reg_1[1029]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2057]),.i2(intermediate_reg_0[2056]),.o(intermediate_reg_1[1028])); 
fsm fsm_inst_1_772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2055]),.i2(intermediate_reg_0[2054]),.o(intermediate_reg_1[1027])); 
mux_module mux_module_inst_1_773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2053]),.i2(intermediate_reg_0[2052]),.o(intermediate_reg_1[1026]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2051]),.i2(intermediate_reg_0[2050]),.o(intermediate_reg_1[1025])); 
fsm fsm_inst_1_775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2049]),.i2(intermediate_reg_0[2048]),.o(intermediate_reg_1[1024])); 
mux_module mux_module_inst_1_776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2047]),.i2(intermediate_reg_0[2046]),.o(intermediate_reg_1[1023]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2045]),.i2(intermediate_reg_0[2044]),.o(intermediate_reg_1[1022]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2043]),.i2(intermediate_reg_0[2042]),.o(intermediate_reg_1[1021]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2041]),.i2(intermediate_reg_0[2040]),.o(intermediate_reg_1[1020]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2039]),.i2(intermediate_reg_0[2038]),.o(intermediate_reg_1[1019])); 
fsm fsm_inst_1_781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2037]),.i2(intermediate_reg_0[2036]),.o(intermediate_reg_1[1018])); 
mux_module mux_module_inst_1_782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2035]),.i2(intermediate_reg_0[2034]),.o(intermediate_reg_1[1017]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2033]),.i2(intermediate_reg_0[2032]),.o(intermediate_reg_1[1016]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2031]),.i2(intermediate_reg_0[2030]),.o(intermediate_reg_1[1015])); 
mux_module mux_module_inst_1_785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2029]),.i2(intermediate_reg_0[2028]),.o(intermediate_reg_1[1014]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2027]),.i2(intermediate_reg_0[2026]),.o(intermediate_reg_1[1013])); 
mux_module mux_module_inst_1_787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2025]),.i2(intermediate_reg_0[2024]),.o(intermediate_reg_1[1012]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2023]),.i2(intermediate_reg_0[2022]),.o(intermediate_reg_1[1011])); 
mux_module mux_module_inst_1_789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2021]),.i2(intermediate_reg_0[2020]),.o(intermediate_reg_1[1010]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2019]),.i2(intermediate_reg_0[2018]),.o(intermediate_reg_1[1009]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2017]),.i2(intermediate_reg_0[2016]),.o(intermediate_reg_1[1008]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2015]),.i2(intermediate_reg_0[2014]),.o(intermediate_reg_1[1007])); 
mux_module mux_module_inst_1_793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2013]),.i2(intermediate_reg_0[2012]),.o(intermediate_reg_1[1006]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2011]),.i2(intermediate_reg_0[2010]),.o(intermediate_reg_1[1005])); 
fsm fsm_inst_1_795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2009]),.i2(intermediate_reg_0[2008]),.o(intermediate_reg_1[1004])); 
mux_module mux_module_inst_1_796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2007]),.i2(intermediate_reg_0[2006]),.o(intermediate_reg_1[1003]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2005]),.i2(intermediate_reg_0[2004]),.o(intermediate_reg_1[1002])); 
mux_module mux_module_inst_1_798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2003]),.i2(intermediate_reg_0[2002]),.o(intermediate_reg_1[1001]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[2001]),.i2(intermediate_reg_0[2000]),.o(intermediate_reg_1[1000])); 
mux_module mux_module_inst_1_800(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1999]),.i2(intermediate_reg_0[1998]),.o(intermediate_reg_1[999]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_801(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1997]),.i2(intermediate_reg_0[1996]),.o(intermediate_reg_1[998])); 
mux_module mux_module_inst_1_802(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1995]),.i2(intermediate_reg_0[1994]),.o(intermediate_reg_1[997]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_803(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1993]),.i2(intermediate_reg_0[1992]),.o(intermediate_reg_1[996])); 
mux_module mux_module_inst_1_804(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1991]),.i2(intermediate_reg_0[1990]),.o(intermediate_reg_1[995]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_805(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1989]),.i2(intermediate_reg_0[1988]),.o(intermediate_reg_1[994]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_806(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1987]),.i2(intermediate_reg_0[1986]),.o(intermediate_reg_1[993]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_807(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1985]),.i2(intermediate_reg_0[1984]),.o(intermediate_reg_1[992])); 
mux_module mux_module_inst_1_808(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1983]),.i2(intermediate_reg_0[1982]),.o(intermediate_reg_1[991]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_809(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1981]),.i2(intermediate_reg_0[1980]),.o(intermediate_reg_1[990]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_810(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1979]),.i2(intermediate_reg_0[1978]),.o(intermediate_reg_1[989])); 
fsm fsm_inst_1_811(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1977]),.i2(intermediate_reg_0[1976]),.o(intermediate_reg_1[988])); 
fsm fsm_inst_1_812(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1975]),.i2(intermediate_reg_0[1974]),.o(intermediate_reg_1[987])); 
mux_module mux_module_inst_1_813(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1973]),.i2(intermediate_reg_0[1972]),.o(intermediate_reg_1[986]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_814(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1971]),.i2(intermediate_reg_0[1970]),.o(intermediate_reg_1[985])); 
mux_module mux_module_inst_1_815(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1969]),.i2(intermediate_reg_0[1968]),.o(intermediate_reg_1[984]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_816(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1967]),.i2(intermediate_reg_0[1966]),.o(intermediate_reg_1[983]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_817(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1965]),.i2(intermediate_reg_0[1964]),.o(intermediate_reg_1[982])); 
fsm fsm_inst_1_818(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1963]),.i2(intermediate_reg_0[1962]),.o(intermediate_reg_1[981])); 
fsm fsm_inst_1_819(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1961]),.i2(intermediate_reg_0[1960]),.o(intermediate_reg_1[980])); 
mux_module mux_module_inst_1_820(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1959]),.i2(intermediate_reg_0[1958]),.o(intermediate_reg_1[979]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_821(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1957]),.i2(intermediate_reg_0[1956]),.o(intermediate_reg_1[978]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_822(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1955]),.i2(intermediate_reg_0[1954]),.o(intermediate_reg_1[977])); 
mux_module mux_module_inst_1_823(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1953]),.i2(intermediate_reg_0[1952]),.o(intermediate_reg_1[976]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_824(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1951]),.i2(intermediate_reg_0[1950]),.o(intermediate_reg_1[975]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_825(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1949]),.i2(intermediate_reg_0[1948]),.o(intermediate_reg_1[974]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_826(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1947]),.i2(intermediate_reg_0[1946]),.o(intermediate_reg_1[973]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_827(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1945]),.i2(intermediate_reg_0[1944]),.o(intermediate_reg_1[972])); 
fsm fsm_inst_1_828(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1943]),.i2(intermediate_reg_0[1942]),.o(intermediate_reg_1[971])); 
mux_module mux_module_inst_1_829(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1941]),.i2(intermediate_reg_0[1940]),.o(intermediate_reg_1[970]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_830(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1939]),.i2(intermediate_reg_0[1938]),.o(intermediate_reg_1[969]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_831(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1937]),.i2(intermediate_reg_0[1936]),.o(intermediate_reg_1[968]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_832(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1935]),.i2(intermediate_reg_0[1934]),.o(intermediate_reg_1[967])); 
mux_module mux_module_inst_1_833(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1933]),.i2(intermediate_reg_0[1932]),.o(intermediate_reg_1[966]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_834(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1931]),.i2(intermediate_reg_0[1930]),.o(intermediate_reg_1[965]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_835(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1929]),.i2(intermediate_reg_0[1928]),.o(intermediate_reg_1[964]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_836(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1927]),.i2(intermediate_reg_0[1926]),.o(intermediate_reg_1[963])); 
fsm fsm_inst_1_837(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1925]),.i2(intermediate_reg_0[1924]),.o(intermediate_reg_1[962])); 
mux_module mux_module_inst_1_838(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1923]),.i2(intermediate_reg_0[1922]),.o(intermediate_reg_1[961]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_839(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1921]),.i2(intermediate_reg_0[1920]),.o(intermediate_reg_1[960]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_840(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1919]),.i2(intermediate_reg_0[1918]),.o(intermediate_reg_1[959]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_841(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1917]),.i2(intermediate_reg_0[1916]),.o(intermediate_reg_1[958])); 
fsm fsm_inst_1_842(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1915]),.i2(intermediate_reg_0[1914]),.o(intermediate_reg_1[957])); 
fsm fsm_inst_1_843(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1913]),.i2(intermediate_reg_0[1912]),.o(intermediate_reg_1[956])); 
mux_module mux_module_inst_1_844(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1911]),.i2(intermediate_reg_0[1910]),.o(intermediate_reg_1[955]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_845(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1909]),.i2(intermediate_reg_0[1908]),.o(intermediate_reg_1[954]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_846(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1907]),.i2(intermediate_reg_0[1906]),.o(intermediate_reg_1[953])); 
mux_module mux_module_inst_1_847(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1905]),.i2(intermediate_reg_0[1904]),.o(intermediate_reg_1[952]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_848(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1903]),.i2(intermediate_reg_0[1902]),.o(intermediate_reg_1[951])); 
mux_module mux_module_inst_1_849(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1901]),.i2(intermediate_reg_0[1900]),.o(intermediate_reg_1[950]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_850(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1899]),.i2(intermediate_reg_0[1898]),.o(intermediate_reg_1[949])); 
mux_module mux_module_inst_1_851(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1897]),.i2(intermediate_reg_0[1896]),.o(intermediate_reg_1[948]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_852(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1895]),.i2(intermediate_reg_0[1894]),.o(intermediate_reg_1[947]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_853(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1893]),.i2(intermediate_reg_0[1892]),.o(intermediate_reg_1[946])); 
fsm fsm_inst_1_854(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1891]),.i2(intermediate_reg_0[1890]),.o(intermediate_reg_1[945])); 
mux_module mux_module_inst_1_855(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1889]),.i2(intermediate_reg_0[1888]),.o(intermediate_reg_1[944]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_856(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1887]),.i2(intermediate_reg_0[1886]),.o(intermediate_reg_1[943])); 
fsm fsm_inst_1_857(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1885]),.i2(intermediate_reg_0[1884]),.o(intermediate_reg_1[942])); 
fsm fsm_inst_1_858(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1883]),.i2(intermediate_reg_0[1882]),.o(intermediate_reg_1[941])); 
mux_module mux_module_inst_1_859(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1881]),.i2(intermediate_reg_0[1880]),.o(intermediate_reg_1[940]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_860(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1879]),.i2(intermediate_reg_0[1878]),.o(intermediate_reg_1[939])); 
fsm fsm_inst_1_861(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1877]),.i2(intermediate_reg_0[1876]),.o(intermediate_reg_1[938])); 
fsm fsm_inst_1_862(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1875]),.i2(intermediate_reg_0[1874]),.o(intermediate_reg_1[937])); 
fsm fsm_inst_1_863(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1873]),.i2(intermediate_reg_0[1872]),.o(intermediate_reg_1[936])); 
mux_module mux_module_inst_1_864(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1871]),.i2(intermediate_reg_0[1870]),.o(intermediate_reg_1[935]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_865(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1869]),.i2(intermediate_reg_0[1868]),.o(intermediate_reg_1[934])); 
fsm fsm_inst_1_866(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1867]),.i2(intermediate_reg_0[1866]),.o(intermediate_reg_1[933])); 
fsm fsm_inst_1_867(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1865]),.i2(intermediate_reg_0[1864]),.o(intermediate_reg_1[932])); 
fsm fsm_inst_1_868(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1863]),.i2(intermediate_reg_0[1862]),.o(intermediate_reg_1[931])); 
mux_module mux_module_inst_1_869(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1861]),.i2(intermediate_reg_0[1860]),.o(intermediate_reg_1[930]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_870(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1859]),.i2(intermediate_reg_0[1858]),.o(intermediate_reg_1[929])); 
mux_module mux_module_inst_1_871(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1857]),.i2(intermediate_reg_0[1856]),.o(intermediate_reg_1[928]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_872(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1855]),.i2(intermediate_reg_0[1854]),.o(intermediate_reg_1[927]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_873(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1853]),.i2(intermediate_reg_0[1852]),.o(intermediate_reg_1[926])); 
mux_module mux_module_inst_1_874(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1851]),.i2(intermediate_reg_0[1850]),.o(intermediate_reg_1[925]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_875(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1849]),.i2(intermediate_reg_0[1848]),.o(intermediate_reg_1[924])); 
mux_module mux_module_inst_1_876(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1847]),.i2(intermediate_reg_0[1846]),.o(intermediate_reg_1[923]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_877(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1845]),.i2(intermediate_reg_0[1844]),.o(intermediate_reg_1[922])); 
mux_module mux_module_inst_1_878(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1843]),.i2(intermediate_reg_0[1842]),.o(intermediate_reg_1[921]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_879(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1841]),.i2(intermediate_reg_0[1840]),.o(intermediate_reg_1[920]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_880(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1839]),.i2(intermediate_reg_0[1838]),.o(intermediate_reg_1[919]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_881(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1837]),.i2(intermediate_reg_0[1836]),.o(intermediate_reg_1[918])); 
fsm fsm_inst_1_882(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1835]),.i2(intermediate_reg_0[1834]),.o(intermediate_reg_1[917])); 
mux_module mux_module_inst_1_883(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1833]),.i2(intermediate_reg_0[1832]),.o(intermediate_reg_1[916]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_884(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1831]),.i2(intermediate_reg_0[1830]),.o(intermediate_reg_1[915])); 
fsm fsm_inst_1_885(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1829]),.i2(intermediate_reg_0[1828]),.o(intermediate_reg_1[914])); 
mux_module mux_module_inst_1_886(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1827]),.i2(intermediate_reg_0[1826]),.o(intermediate_reg_1[913]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_887(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1825]),.i2(intermediate_reg_0[1824]),.o(intermediate_reg_1[912])); 
mux_module mux_module_inst_1_888(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1823]),.i2(intermediate_reg_0[1822]),.o(intermediate_reg_1[911]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_889(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1821]),.i2(intermediate_reg_0[1820]),.o(intermediate_reg_1[910]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_890(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1819]),.i2(intermediate_reg_0[1818]),.o(intermediate_reg_1[909]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_891(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1817]),.i2(intermediate_reg_0[1816]),.o(intermediate_reg_1[908])); 
fsm fsm_inst_1_892(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1815]),.i2(intermediate_reg_0[1814]),.o(intermediate_reg_1[907])); 
mux_module mux_module_inst_1_893(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1813]),.i2(intermediate_reg_0[1812]),.o(intermediate_reg_1[906]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_894(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1811]),.i2(intermediate_reg_0[1810]),.o(intermediate_reg_1[905]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_895(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1809]),.i2(intermediate_reg_0[1808]),.o(intermediate_reg_1[904])); 
fsm fsm_inst_1_896(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1807]),.i2(intermediate_reg_0[1806]),.o(intermediate_reg_1[903])); 
mux_module mux_module_inst_1_897(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1805]),.i2(intermediate_reg_0[1804]),.o(intermediate_reg_1[902]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_898(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1803]),.i2(intermediate_reg_0[1802]),.o(intermediate_reg_1[901])); 
mux_module mux_module_inst_1_899(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1801]),.i2(intermediate_reg_0[1800]),.o(intermediate_reg_1[900]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_900(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1799]),.i2(intermediate_reg_0[1798]),.o(intermediate_reg_1[899])); 
fsm fsm_inst_1_901(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1797]),.i2(intermediate_reg_0[1796]),.o(intermediate_reg_1[898])); 
fsm fsm_inst_1_902(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1795]),.i2(intermediate_reg_0[1794]),.o(intermediate_reg_1[897])); 
mux_module mux_module_inst_1_903(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1793]),.i2(intermediate_reg_0[1792]),.o(intermediate_reg_1[896]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_904(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1791]),.i2(intermediate_reg_0[1790]),.o(intermediate_reg_1[895]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_905(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1789]),.i2(intermediate_reg_0[1788]),.o(intermediate_reg_1[894]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_906(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1787]),.i2(intermediate_reg_0[1786]),.o(intermediate_reg_1[893])); 
fsm fsm_inst_1_907(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1785]),.i2(intermediate_reg_0[1784]),.o(intermediate_reg_1[892])); 
mux_module mux_module_inst_1_908(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1783]),.i2(intermediate_reg_0[1782]),.o(intermediate_reg_1[891]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_909(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1781]),.i2(intermediate_reg_0[1780]),.o(intermediate_reg_1[890])); 
fsm fsm_inst_1_910(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1779]),.i2(intermediate_reg_0[1778]),.o(intermediate_reg_1[889])); 
mux_module mux_module_inst_1_911(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1777]),.i2(intermediate_reg_0[1776]),.o(intermediate_reg_1[888]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_912(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1775]),.i2(intermediate_reg_0[1774]),.o(intermediate_reg_1[887]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_913(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1773]),.i2(intermediate_reg_0[1772]),.o(intermediate_reg_1[886])); 
fsm fsm_inst_1_914(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1771]),.i2(intermediate_reg_0[1770]),.o(intermediate_reg_1[885])); 
fsm fsm_inst_1_915(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1769]),.i2(intermediate_reg_0[1768]),.o(intermediate_reg_1[884])); 
mux_module mux_module_inst_1_916(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1767]),.i2(intermediate_reg_0[1766]),.o(intermediate_reg_1[883]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_917(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1765]),.i2(intermediate_reg_0[1764]),.o(intermediate_reg_1[882]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_918(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1763]),.i2(intermediate_reg_0[1762]),.o(intermediate_reg_1[881])); 
fsm fsm_inst_1_919(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1761]),.i2(intermediate_reg_0[1760]),.o(intermediate_reg_1[880])); 
fsm fsm_inst_1_920(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1759]),.i2(intermediate_reg_0[1758]),.o(intermediate_reg_1[879])); 
fsm fsm_inst_1_921(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1757]),.i2(intermediate_reg_0[1756]),.o(intermediate_reg_1[878])); 
mux_module mux_module_inst_1_922(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1755]),.i2(intermediate_reg_0[1754]),.o(intermediate_reg_1[877]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_923(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1753]),.i2(intermediate_reg_0[1752]),.o(intermediate_reg_1[876]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_924(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1751]),.i2(intermediate_reg_0[1750]),.o(intermediate_reg_1[875])); 
fsm fsm_inst_1_925(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1749]),.i2(intermediate_reg_0[1748]),.o(intermediate_reg_1[874])); 
mux_module mux_module_inst_1_926(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1747]),.i2(intermediate_reg_0[1746]),.o(intermediate_reg_1[873]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_927(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1745]),.i2(intermediate_reg_0[1744]),.o(intermediate_reg_1[872]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_928(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1743]),.i2(intermediate_reg_0[1742]),.o(intermediate_reg_1[871]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_929(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1741]),.i2(intermediate_reg_0[1740]),.o(intermediate_reg_1[870]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_930(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1739]),.i2(intermediate_reg_0[1738]),.o(intermediate_reg_1[869])); 
fsm fsm_inst_1_931(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1737]),.i2(intermediate_reg_0[1736]),.o(intermediate_reg_1[868])); 
fsm fsm_inst_1_932(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1735]),.i2(intermediate_reg_0[1734]),.o(intermediate_reg_1[867])); 
fsm fsm_inst_1_933(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1733]),.i2(intermediate_reg_0[1732]),.o(intermediate_reg_1[866])); 
mux_module mux_module_inst_1_934(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1731]),.i2(intermediate_reg_0[1730]),.o(intermediate_reg_1[865]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_935(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1729]),.i2(intermediate_reg_0[1728]),.o(intermediate_reg_1[864])); 
mux_module mux_module_inst_1_936(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1727]),.i2(intermediate_reg_0[1726]),.o(intermediate_reg_1[863]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_937(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1725]),.i2(intermediate_reg_0[1724]),.o(intermediate_reg_1[862])); 
fsm fsm_inst_1_938(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1723]),.i2(intermediate_reg_0[1722]),.o(intermediate_reg_1[861])); 
mux_module mux_module_inst_1_939(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1721]),.i2(intermediate_reg_0[1720]),.o(intermediate_reg_1[860]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_940(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1719]),.i2(intermediate_reg_0[1718]),.o(intermediate_reg_1[859]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_941(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1717]),.i2(intermediate_reg_0[1716]),.o(intermediate_reg_1[858]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_942(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1715]),.i2(intermediate_reg_0[1714]),.o(intermediate_reg_1[857]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_943(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1713]),.i2(intermediate_reg_0[1712]),.o(intermediate_reg_1[856])); 
fsm fsm_inst_1_944(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1711]),.i2(intermediate_reg_0[1710]),.o(intermediate_reg_1[855])); 
fsm fsm_inst_1_945(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1709]),.i2(intermediate_reg_0[1708]),.o(intermediate_reg_1[854])); 
mux_module mux_module_inst_1_946(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1707]),.i2(intermediate_reg_0[1706]),.o(intermediate_reg_1[853]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_947(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1705]),.i2(intermediate_reg_0[1704]),.o(intermediate_reg_1[852]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_948(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1703]),.i2(intermediate_reg_0[1702]),.o(intermediate_reg_1[851]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_949(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1701]),.i2(intermediate_reg_0[1700]),.o(intermediate_reg_1[850]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_950(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1699]),.i2(intermediate_reg_0[1698]),.o(intermediate_reg_1[849]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_951(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1697]),.i2(intermediate_reg_0[1696]),.o(intermediate_reg_1[848])); 
fsm fsm_inst_1_952(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1695]),.i2(intermediate_reg_0[1694]),.o(intermediate_reg_1[847])); 
fsm fsm_inst_1_953(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1693]),.i2(intermediate_reg_0[1692]),.o(intermediate_reg_1[846])); 
fsm fsm_inst_1_954(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1691]),.i2(intermediate_reg_0[1690]),.o(intermediate_reg_1[845])); 
mux_module mux_module_inst_1_955(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1689]),.i2(intermediate_reg_0[1688]),.o(intermediate_reg_1[844]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_956(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1687]),.i2(intermediate_reg_0[1686]),.o(intermediate_reg_1[843])); 
mux_module mux_module_inst_1_957(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1685]),.i2(intermediate_reg_0[1684]),.o(intermediate_reg_1[842]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_958(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1683]),.i2(intermediate_reg_0[1682]),.o(intermediate_reg_1[841])); 
fsm fsm_inst_1_959(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1681]),.i2(intermediate_reg_0[1680]),.o(intermediate_reg_1[840])); 
mux_module mux_module_inst_1_960(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1679]),.i2(intermediate_reg_0[1678]),.o(intermediate_reg_1[839]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_961(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1677]),.i2(intermediate_reg_0[1676]),.o(intermediate_reg_1[838])); 
mux_module mux_module_inst_1_962(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1675]),.i2(intermediate_reg_0[1674]),.o(intermediate_reg_1[837]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_963(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1673]),.i2(intermediate_reg_0[1672]),.o(intermediate_reg_1[836])); 
mux_module mux_module_inst_1_964(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1671]),.i2(intermediate_reg_0[1670]),.o(intermediate_reg_1[835]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_965(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1669]),.i2(intermediate_reg_0[1668]),.o(intermediate_reg_1[834])); 
mux_module mux_module_inst_1_966(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1667]),.i2(intermediate_reg_0[1666]),.o(intermediate_reg_1[833]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_967(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1665]),.i2(intermediate_reg_0[1664]),.o(intermediate_reg_1[832]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_968(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1663]),.i2(intermediate_reg_0[1662]),.o(intermediate_reg_1[831])); 
mux_module mux_module_inst_1_969(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1661]),.i2(intermediate_reg_0[1660]),.o(intermediate_reg_1[830]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_970(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1659]),.i2(intermediate_reg_0[1658]),.o(intermediate_reg_1[829]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_971(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1657]),.i2(intermediate_reg_0[1656]),.o(intermediate_reg_1[828]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_972(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1655]),.i2(intermediate_reg_0[1654]),.o(intermediate_reg_1[827]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_973(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1653]),.i2(intermediate_reg_0[1652]),.o(intermediate_reg_1[826])); 
fsm fsm_inst_1_974(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1651]),.i2(intermediate_reg_0[1650]),.o(intermediate_reg_1[825])); 
mux_module mux_module_inst_1_975(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1649]),.i2(intermediate_reg_0[1648]),.o(intermediate_reg_1[824]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_976(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1647]),.i2(intermediate_reg_0[1646]),.o(intermediate_reg_1[823])); 
fsm fsm_inst_1_977(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1645]),.i2(intermediate_reg_0[1644]),.o(intermediate_reg_1[822])); 
fsm fsm_inst_1_978(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1643]),.i2(intermediate_reg_0[1642]),.o(intermediate_reg_1[821])); 
fsm fsm_inst_1_979(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1641]),.i2(intermediate_reg_0[1640]),.o(intermediate_reg_1[820])); 
fsm fsm_inst_1_980(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1639]),.i2(intermediate_reg_0[1638]),.o(intermediate_reg_1[819])); 
mux_module mux_module_inst_1_981(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1637]),.i2(intermediate_reg_0[1636]),.o(intermediate_reg_1[818]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_982(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1635]),.i2(intermediate_reg_0[1634]),.o(intermediate_reg_1[817])); 
mux_module mux_module_inst_1_983(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1633]),.i2(intermediate_reg_0[1632]),.o(intermediate_reg_1[816]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_984(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1631]),.i2(intermediate_reg_0[1630]),.o(intermediate_reg_1[815]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_985(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1629]),.i2(intermediate_reg_0[1628]),.o(intermediate_reg_1[814]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_986(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1627]),.i2(intermediate_reg_0[1626]),.o(intermediate_reg_1[813]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_987(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1625]),.i2(intermediate_reg_0[1624]),.o(intermediate_reg_1[812]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_988(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1623]),.i2(intermediate_reg_0[1622]),.o(intermediate_reg_1[811]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_989(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1621]),.i2(intermediate_reg_0[1620]),.o(intermediate_reg_1[810])); 
fsm fsm_inst_1_990(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1619]),.i2(intermediate_reg_0[1618]),.o(intermediate_reg_1[809])); 
fsm fsm_inst_1_991(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1617]),.i2(intermediate_reg_0[1616]),.o(intermediate_reg_1[808])); 
fsm fsm_inst_1_992(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1615]),.i2(intermediate_reg_0[1614]),.o(intermediate_reg_1[807])); 
mux_module mux_module_inst_1_993(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1613]),.i2(intermediate_reg_0[1612]),.o(intermediate_reg_1[806]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_994(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1611]),.i2(intermediate_reg_0[1610]),.o(intermediate_reg_1[805])); 
mux_module mux_module_inst_1_995(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1609]),.i2(intermediate_reg_0[1608]),.o(intermediate_reg_1[804]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_996(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1607]),.i2(intermediate_reg_0[1606]),.o(intermediate_reg_1[803]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_997(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1605]),.i2(intermediate_reg_0[1604]),.o(intermediate_reg_1[802]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_998(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1603]),.i2(intermediate_reg_0[1602]),.o(intermediate_reg_1[801])); 
mux_module mux_module_inst_1_999(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1601]),.i2(intermediate_reg_0[1600]),.o(intermediate_reg_1[800]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1000(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1599]),.i2(intermediate_reg_0[1598]),.o(intermediate_reg_1[799]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1001(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1597]),.i2(intermediate_reg_0[1596]),.o(intermediate_reg_1[798])); 
fsm fsm_inst_1_1002(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1595]),.i2(intermediate_reg_0[1594]),.o(intermediate_reg_1[797])); 
mux_module mux_module_inst_1_1003(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1593]),.i2(intermediate_reg_0[1592]),.o(intermediate_reg_1[796]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1004(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1591]),.i2(intermediate_reg_0[1590]),.o(intermediate_reg_1[795])); 
mux_module mux_module_inst_1_1005(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1589]),.i2(intermediate_reg_0[1588]),.o(intermediate_reg_1[794]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1006(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1587]),.i2(intermediate_reg_0[1586]),.o(intermediate_reg_1[793])); 
mux_module mux_module_inst_1_1007(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1585]),.i2(intermediate_reg_0[1584]),.o(intermediate_reg_1[792]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1008(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1583]),.i2(intermediate_reg_0[1582]),.o(intermediate_reg_1[791]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1009(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1581]),.i2(intermediate_reg_0[1580]),.o(intermediate_reg_1[790]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1010(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1579]),.i2(intermediate_reg_0[1578]),.o(intermediate_reg_1[789])); 
fsm fsm_inst_1_1011(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1577]),.i2(intermediate_reg_0[1576]),.o(intermediate_reg_1[788])); 
fsm fsm_inst_1_1012(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1575]),.i2(intermediate_reg_0[1574]),.o(intermediate_reg_1[787])); 
fsm fsm_inst_1_1013(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1573]),.i2(intermediate_reg_0[1572]),.o(intermediate_reg_1[786])); 
fsm fsm_inst_1_1014(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1571]),.i2(intermediate_reg_0[1570]),.o(intermediate_reg_1[785])); 
mux_module mux_module_inst_1_1015(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1569]),.i2(intermediate_reg_0[1568]),.o(intermediate_reg_1[784]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1016(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1567]),.i2(intermediate_reg_0[1566]),.o(intermediate_reg_1[783])); 
fsm fsm_inst_1_1017(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1565]),.i2(intermediate_reg_0[1564]),.o(intermediate_reg_1[782])); 
fsm fsm_inst_1_1018(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1563]),.i2(intermediate_reg_0[1562]),.o(intermediate_reg_1[781])); 
fsm fsm_inst_1_1019(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1561]),.i2(intermediate_reg_0[1560]),.o(intermediate_reg_1[780])); 
fsm fsm_inst_1_1020(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1559]),.i2(intermediate_reg_0[1558]),.o(intermediate_reg_1[779])); 
mux_module mux_module_inst_1_1021(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1557]),.i2(intermediate_reg_0[1556]),.o(intermediate_reg_1[778]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1022(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1555]),.i2(intermediate_reg_0[1554]),.o(intermediate_reg_1[777])); 
fsm fsm_inst_1_1023(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1553]),.i2(intermediate_reg_0[1552]),.o(intermediate_reg_1[776])); 
fsm fsm_inst_1_1024(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1551]),.i2(intermediate_reg_0[1550]),.o(intermediate_reg_1[775])); 
fsm fsm_inst_1_1025(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1549]),.i2(intermediate_reg_0[1548]),.o(intermediate_reg_1[774])); 
mux_module mux_module_inst_1_1026(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1547]),.i2(intermediate_reg_0[1546]),.o(intermediate_reg_1[773]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1027(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1545]),.i2(intermediate_reg_0[1544]),.o(intermediate_reg_1[772])); 
fsm fsm_inst_1_1028(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1543]),.i2(intermediate_reg_0[1542]),.o(intermediate_reg_1[771])); 
mux_module mux_module_inst_1_1029(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1541]),.i2(intermediate_reg_0[1540]),.o(intermediate_reg_1[770]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1030(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1539]),.i2(intermediate_reg_0[1538]),.o(intermediate_reg_1[769]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1031(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1537]),.i2(intermediate_reg_0[1536]),.o(intermediate_reg_1[768]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1032(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1535]),.i2(intermediate_reg_0[1534]),.o(intermediate_reg_1[767]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1033(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1533]),.i2(intermediate_reg_0[1532]),.o(intermediate_reg_1[766])); 
fsm fsm_inst_1_1034(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1531]),.i2(intermediate_reg_0[1530]),.o(intermediate_reg_1[765])); 
fsm fsm_inst_1_1035(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1529]),.i2(intermediate_reg_0[1528]),.o(intermediate_reg_1[764])); 
fsm fsm_inst_1_1036(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1527]),.i2(intermediate_reg_0[1526]),.o(intermediate_reg_1[763])); 
fsm fsm_inst_1_1037(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1525]),.i2(intermediate_reg_0[1524]),.o(intermediate_reg_1[762])); 
mux_module mux_module_inst_1_1038(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1523]),.i2(intermediate_reg_0[1522]),.o(intermediate_reg_1[761]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1039(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1521]),.i2(intermediate_reg_0[1520]),.o(intermediate_reg_1[760])); 
fsm fsm_inst_1_1040(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1519]),.i2(intermediate_reg_0[1518]),.o(intermediate_reg_1[759])); 
mux_module mux_module_inst_1_1041(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1517]),.i2(intermediate_reg_0[1516]),.o(intermediate_reg_1[758]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1042(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1515]),.i2(intermediate_reg_0[1514]),.o(intermediate_reg_1[757]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1043(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1513]),.i2(intermediate_reg_0[1512]),.o(intermediate_reg_1[756])); 
mux_module mux_module_inst_1_1044(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1511]),.i2(intermediate_reg_0[1510]),.o(intermediate_reg_1[755]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1045(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1509]),.i2(intermediate_reg_0[1508]),.o(intermediate_reg_1[754]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1046(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1507]),.i2(intermediate_reg_0[1506]),.o(intermediate_reg_1[753]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1047(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1505]),.i2(intermediate_reg_0[1504]),.o(intermediate_reg_1[752])); 
mux_module mux_module_inst_1_1048(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1503]),.i2(intermediate_reg_0[1502]),.o(intermediate_reg_1[751]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1049(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1501]),.i2(intermediate_reg_0[1500]),.o(intermediate_reg_1[750])); 
fsm fsm_inst_1_1050(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1499]),.i2(intermediate_reg_0[1498]),.o(intermediate_reg_1[749])); 
fsm fsm_inst_1_1051(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1497]),.i2(intermediate_reg_0[1496]),.o(intermediate_reg_1[748])); 
mux_module mux_module_inst_1_1052(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1495]),.i2(intermediate_reg_0[1494]),.o(intermediate_reg_1[747]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1053(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1493]),.i2(intermediate_reg_0[1492]),.o(intermediate_reg_1[746]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1054(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1491]),.i2(intermediate_reg_0[1490]),.o(intermediate_reg_1[745]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1055(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1489]),.i2(intermediate_reg_0[1488]),.o(intermediate_reg_1[744])); 
mux_module mux_module_inst_1_1056(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1487]),.i2(intermediate_reg_0[1486]),.o(intermediate_reg_1[743]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1057(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1485]),.i2(intermediate_reg_0[1484]),.o(intermediate_reg_1[742])); 
fsm fsm_inst_1_1058(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1483]),.i2(intermediate_reg_0[1482]),.o(intermediate_reg_1[741])); 
mux_module mux_module_inst_1_1059(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1481]),.i2(intermediate_reg_0[1480]),.o(intermediate_reg_1[740]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1060(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1479]),.i2(intermediate_reg_0[1478]),.o(intermediate_reg_1[739]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1061(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1477]),.i2(intermediate_reg_0[1476]),.o(intermediate_reg_1[738]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1062(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1475]),.i2(intermediate_reg_0[1474]),.o(intermediate_reg_1[737]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1063(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1473]),.i2(intermediate_reg_0[1472]),.o(intermediate_reg_1[736]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1064(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1471]),.i2(intermediate_reg_0[1470]),.o(intermediate_reg_1[735]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1065(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1469]),.i2(intermediate_reg_0[1468]),.o(intermediate_reg_1[734])); 
mux_module mux_module_inst_1_1066(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1467]),.i2(intermediate_reg_0[1466]),.o(intermediate_reg_1[733]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1067(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1465]),.i2(intermediate_reg_0[1464]),.o(intermediate_reg_1[732]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1068(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1463]),.i2(intermediate_reg_0[1462]),.o(intermediate_reg_1[731])); 
fsm fsm_inst_1_1069(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1461]),.i2(intermediate_reg_0[1460]),.o(intermediate_reg_1[730])); 
mux_module mux_module_inst_1_1070(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1459]),.i2(intermediate_reg_0[1458]),.o(intermediate_reg_1[729]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1071(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1457]),.i2(intermediate_reg_0[1456]),.o(intermediate_reg_1[728]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1072(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1455]),.i2(intermediate_reg_0[1454]),.o(intermediate_reg_1[727]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1073(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1453]),.i2(intermediate_reg_0[1452]),.o(intermediate_reg_1[726])); 
mux_module mux_module_inst_1_1074(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1451]),.i2(intermediate_reg_0[1450]),.o(intermediate_reg_1[725]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1075(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1449]),.i2(intermediate_reg_0[1448]),.o(intermediate_reg_1[724]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1076(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1447]),.i2(intermediate_reg_0[1446]),.o(intermediate_reg_1[723])); 
fsm fsm_inst_1_1077(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1445]),.i2(intermediate_reg_0[1444]),.o(intermediate_reg_1[722])); 
mux_module mux_module_inst_1_1078(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1443]),.i2(intermediate_reg_0[1442]),.o(intermediate_reg_1[721]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1079(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1441]),.i2(intermediate_reg_0[1440]),.o(intermediate_reg_1[720]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1080(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1439]),.i2(intermediate_reg_0[1438]),.o(intermediate_reg_1[719])); 
mux_module mux_module_inst_1_1081(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1437]),.i2(intermediate_reg_0[1436]),.o(intermediate_reg_1[718]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1082(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1435]),.i2(intermediate_reg_0[1434]),.o(intermediate_reg_1[717])); 
mux_module mux_module_inst_1_1083(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1433]),.i2(intermediate_reg_0[1432]),.o(intermediate_reg_1[716]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1084(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1431]),.i2(intermediate_reg_0[1430]),.o(intermediate_reg_1[715])); 
mux_module mux_module_inst_1_1085(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1429]),.i2(intermediate_reg_0[1428]),.o(intermediate_reg_1[714]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1086(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1427]),.i2(intermediate_reg_0[1426]),.o(intermediate_reg_1[713])); 
fsm fsm_inst_1_1087(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1425]),.i2(intermediate_reg_0[1424]),.o(intermediate_reg_1[712])); 
fsm fsm_inst_1_1088(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1423]),.i2(intermediate_reg_0[1422]),.o(intermediate_reg_1[711])); 
fsm fsm_inst_1_1089(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1421]),.i2(intermediate_reg_0[1420]),.o(intermediate_reg_1[710])); 
mux_module mux_module_inst_1_1090(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1419]),.i2(intermediate_reg_0[1418]),.o(intermediate_reg_1[709]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1091(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1417]),.i2(intermediate_reg_0[1416]),.o(intermediate_reg_1[708])); 
fsm fsm_inst_1_1092(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1415]),.i2(intermediate_reg_0[1414]),.o(intermediate_reg_1[707])); 
mux_module mux_module_inst_1_1093(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1413]),.i2(intermediate_reg_0[1412]),.o(intermediate_reg_1[706]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1094(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1411]),.i2(intermediate_reg_0[1410]),.o(intermediate_reg_1[705])); 
mux_module mux_module_inst_1_1095(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1409]),.i2(intermediate_reg_0[1408]),.o(intermediate_reg_1[704]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1096(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1407]),.i2(intermediate_reg_0[1406]),.o(intermediate_reg_1[703])); 
fsm fsm_inst_1_1097(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1405]),.i2(intermediate_reg_0[1404]),.o(intermediate_reg_1[702])); 
fsm fsm_inst_1_1098(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1403]),.i2(intermediate_reg_0[1402]),.o(intermediate_reg_1[701])); 
mux_module mux_module_inst_1_1099(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1401]),.i2(intermediate_reg_0[1400]),.o(intermediate_reg_1[700]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1100(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1399]),.i2(intermediate_reg_0[1398]),.o(intermediate_reg_1[699])); 
mux_module mux_module_inst_1_1101(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1397]),.i2(intermediate_reg_0[1396]),.o(intermediate_reg_1[698]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1102(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1395]),.i2(intermediate_reg_0[1394]),.o(intermediate_reg_1[697]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1103(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1393]),.i2(intermediate_reg_0[1392]),.o(intermediate_reg_1[696])); 
mux_module mux_module_inst_1_1104(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1391]),.i2(intermediate_reg_0[1390]),.o(intermediate_reg_1[695]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1105(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1389]),.i2(intermediate_reg_0[1388]),.o(intermediate_reg_1[694])); 
fsm fsm_inst_1_1106(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1387]),.i2(intermediate_reg_0[1386]),.o(intermediate_reg_1[693])); 
fsm fsm_inst_1_1107(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1385]),.i2(intermediate_reg_0[1384]),.o(intermediate_reg_1[692])); 
fsm fsm_inst_1_1108(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1383]),.i2(intermediate_reg_0[1382]),.o(intermediate_reg_1[691])); 
fsm fsm_inst_1_1109(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1381]),.i2(intermediate_reg_0[1380]),.o(intermediate_reg_1[690])); 
fsm fsm_inst_1_1110(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1379]),.i2(intermediate_reg_0[1378]),.o(intermediate_reg_1[689])); 
mux_module mux_module_inst_1_1111(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1377]),.i2(intermediate_reg_0[1376]),.o(intermediate_reg_1[688]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1112(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1375]),.i2(intermediate_reg_0[1374]),.o(intermediate_reg_1[687]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1113(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1373]),.i2(intermediate_reg_0[1372]),.o(intermediate_reg_1[686]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1114(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1371]),.i2(intermediate_reg_0[1370]),.o(intermediate_reg_1[685])); 
mux_module mux_module_inst_1_1115(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1369]),.i2(intermediate_reg_0[1368]),.o(intermediate_reg_1[684]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1116(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1367]),.i2(intermediate_reg_0[1366]),.o(intermediate_reg_1[683]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1117(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1365]),.i2(intermediate_reg_0[1364]),.o(intermediate_reg_1[682]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1118(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1363]),.i2(intermediate_reg_0[1362]),.o(intermediate_reg_1[681])); 
fsm fsm_inst_1_1119(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1361]),.i2(intermediate_reg_0[1360]),.o(intermediate_reg_1[680])); 
fsm fsm_inst_1_1120(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1359]),.i2(intermediate_reg_0[1358]),.o(intermediate_reg_1[679])); 
fsm fsm_inst_1_1121(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1357]),.i2(intermediate_reg_0[1356]),.o(intermediate_reg_1[678])); 
mux_module mux_module_inst_1_1122(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1355]),.i2(intermediate_reg_0[1354]),.o(intermediate_reg_1[677]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1123(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1353]),.i2(intermediate_reg_0[1352]),.o(intermediate_reg_1[676]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1124(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1351]),.i2(intermediate_reg_0[1350]),.o(intermediate_reg_1[675]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1125(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1349]),.i2(intermediate_reg_0[1348]),.o(intermediate_reg_1[674])); 
fsm fsm_inst_1_1126(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1347]),.i2(intermediate_reg_0[1346]),.o(intermediate_reg_1[673])); 
fsm fsm_inst_1_1127(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1345]),.i2(intermediate_reg_0[1344]),.o(intermediate_reg_1[672])); 
mux_module mux_module_inst_1_1128(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1343]),.i2(intermediate_reg_0[1342]),.o(intermediate_reg_1[671]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1129(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1341]),.i2(intermediate_reg_0[1340]),.o(intermediate_reg_1[670]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1130(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1339]),.i2(intermediate_reg_0[1338]),.o(intermediate_reg_1[669]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1131(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1337]),.i2(intermediate_reg_0[1336]),.o(intermediate_reg_1[668])); 
fsm fsm_inst_1_1132(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1335]),.i2(intermediate_reg_0[1334]),.o(intermediate_reg_1[667])); 
mux_module mux_module_inst_1_1133(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1333]),.i2(intermediate_reg_0[1332]),.o(intermediate_reg_1[666]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1134(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1331]),.i2(intermediate_reg_0[1330]),.o(intermediate_reg_1[665]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1135(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1329]),.i2(intermediate_reg_0[1328]),.o(intermediate_reg_1[664]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1136(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1327]),.i2(intermediate_reg_0[1326]),.o(intermediate_reg_1[663])); 
fsm fsm_inst_1_1137(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1325]),.i2(intermediate_reg_0[1324]),.o(intermediate_reg_1[662])); 
mux_module mux_module_inst_1_1138(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1323]),.i2(intermediate_reg_0[1322]),.o(intermediate_reg_1[661]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1139(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1321]),.i2(intermediate_reg_0[1320]),.o(intermediate_reg_1[660])); 
fsm fsm_inst_1_1140(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1319]),.i2(intermediate_reg_0[1318]),.o(intermediate_reg_1[659])); 
fsm fsm_inst_1_1141(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1317]),.i2(intermediate_reg_0[1316]),.o(intermediate_reg_1[658])); 
mux_module mux_module_inst_1_1142(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1315]),.i2(intermediate_reg_0[1314]),.o(intermediate_reg_1[657]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1143(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1313]),.i2(intermediate_reg_0[1312]),.o(intermediate_reg_1[656])); 
fsm fsm_inst_1_1144(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1311]),.i2(intermediate_reg_0[1310]),.o(intermediate_reg_1[655])); 
mux_module mux_module_inst_1_1145(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1309]),.i2(intermediate_reg_0[1308]),.o(intermediate_reg_1[654]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1146(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1307]),.i2(intermediate_reg_0[1306]),.o(intermediate_reg_1[653]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1147(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1305]),.i2(intermediate_reg_0[1304]),.o(intermediate_reg_1[652])); 
mux_module mux_module_inst_1_1148(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1303]),.i2(intermediate_reg_0[1302]),.o(intermediate_reg_1[651]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1149(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1301]),.i2(intermediate_reg_0[1300]),.o(intermediate_reg_1[650]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1150(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1299]),.i2(intermediate_reg_0[1298]),.o(intermediate_reg_1[649]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1151(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1297]),.i2(intermediate_reg_0[1296]),.o(intermediate_reg_1[648]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1152(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1295]),.i2(intermediate_reg_0[1294]),.o(intermediate_reg_1[647])); 
mux_module mux_module_inst_1_1153(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1293]),.i2(intermediate_reg_0[1292]),.o(intermediate_reg_1[646]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1154(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1291]),.i2(intermediate_reg_0[1290]),.o(intermediate_reg_1[645]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1155(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1289]),.i2(intermediate_reg_0[1288]),.o(intermediate_reg_1[644])); 
fsm fsm_inst_1_1156(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1287]),.i2(intermediate_reg_0[1286]),.o(intermediate_reg_1[643])); 
mux_module mux_module_inst_1_1157(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1285]),.i2(intermediate_reg_0[1284]),.o(intermediate_reg_1[642]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1158(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1283]),.i2(intermediate_reg_0[1282]),.o(intermediate_reg_1[641])); 
mux_module mux_module_inst_1_1159(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1281]),.i2(intermediate_reg_0[1280]),.o(intermediate_reg_1[640]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1160(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1279]),.i2(intermediate_reg_0[1278]),.o(intermediate_reg_1[639])); 
mux_module mux_module_inst_1_1161(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1277]),.i2(intermediate_reg_0[1276]),.o(intermediate_reg_1[638]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1162(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1275]),.i2(intermediate_reg_0[1274]),.o(intermediate_reg_1[637])); 
mux_module mux_module_inst_1_1163(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1273]),.i2(intermediate_reg_0[1272]),.o(intermediate_reg_1[636]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1164(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1271]),.i2(intermediate_reg_0[1270]),.o(intermediate_reg_1[635]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1165(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1269]),.i2(intermediate_reg_0[1268]),.o(intermediate_reg_1[634]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1166(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1267]),.i2(intermediate_reg_0[1266]),.o(intermediate_reg_1[633]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1167(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1265]),.i2(intermediate_reg_0[1264]),.o(intermediate_reg_1[632]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1168(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1263]),.i2(intermediate_reg_0[1262]),.o(intermediate_reg_1[631])); 
fsm fsm_inst_1_1169(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1261]),.i2(intermediate_reg_0[1260]),.o(intermediate_reg_1[630])); 
mux_module mux_module_inst_1_1170(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1259]),.i2(intermediate_reg_0[1258]),.o(intermediate_reg_1[629]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1171(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1257]),.i2(intermediate_reg_0[1256]),.o(intermediate_reg_1[628]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1172(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1255]),.i2(intermediate_reg_0[1254]),.o(intermediate_reg_1[627])); 
mux_module mux_module_inst_1_1173(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1253]),.i2(intermediate_reg_0[1252]),.o(intermediate_reg_1[626]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1174(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1251]),.i2(intermediate_reg_0[1250]),.o(intermediate_reg_1[625])); 
fsm fsm_inst_1_1175(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1249]),.i2(intermediate_reg_0[1248]),.o(intermediate_reg_1[624])); 
fsm fsm_inst_1_1176(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1247]),.i2(intermediate_reg_0[1246]),.o(intermediate_reg_1[623])); 
fsm fsm_inst_1_1177(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1245]),.i2(intermediate_reg_0[1244]),.o(intermediate_reg_1[622])); 
mux_module mux_module_inst_1_1178(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1243]),.i2(intermediate_reg_0[1242]),.o(intermediate_reg_1[621]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1179(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1241]),.i2(intermediate_reg_0[1240]),.o(intermediate_reg_1[620]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1180(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1239]),.i2(intermediate_reg_0[1238]),.o(intermediate_reg_1[619])); 
fsm fsm_inst_1_1181(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1237]),.i2(intermediate_reg_0[1236]),.o(intermediate_reg_1[618])); 
fsm fsm_inst_1_1182(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1235]),.i2(intermediate_reg_0[1234]),.o(intermediate_reg_1[617])); 
fsm fsm_inst_1_1183(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1233]),.i2(intermediate_reg_0[1232]),.o(intermediate_reg_1[616])); 
mux_module mux_module_inst_1_1184(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1231]),.i2(intermediate_reg_0[1230]),.o(intermediate_reg_1[615]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1185(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1229]),.i2(intermediate_reg_0[1228]),.o(intermediate_reg_1[614])); 
fsm fsm_inst_1_1186(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1227]),.i2(intermediate_reg_0[1226]),.o(intermediate_reg_1[613])); 
mux_module mux_module_inst_1_1187(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1225]),.i2(intermediate_reg_0[1224]),.o(intermediate_reg_1[612]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1188(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1223]),.i2(intermediate_reg_0[1222]),.o(intermediate_reg_1[611])); 
fsm fsm_inst_1_1189(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1221]),.i2(intermediate_reg_0[1220]),.o(intermediate_reg_1[610])); 
mux_module mux_module_inst_1_1190(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1219]),.i2(intermediate_reg_0[1218]),.o(intermediate_reg_1[609]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1191(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1217]),.i2(intermediate_reg_0[1216]),.o(intermediate_reg_1[608])); 
fsm fsm_inst_1_1192(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1215]),.i2(intermediate_reg_0[1214]),.o(intermediate_reg_1[607])); 
mux_module mux_module_inst_1_1193(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1213]),.i2(intermediate_reg_0[1212]),.o(intermediate_reg_1[606]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1194(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1211]),.i2(intermediate_reg_0[1210]),.o(intermediate_reg_1[605]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1195(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1209]),.i2(intermediate_reg_0[1208]),.o(intermediate_reg_1[604]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1196(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1207]),.i2(intermediate_reg_0[1206]),.o(intermediate_reg_1[603]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1197(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1205]),.i2(intermediate_reg_0[1204]),.o(intermediate_reg_1[602]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1198(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1203]),.i2(intermediate_reg_0[1202]),.o(intermediate_reg_1[601])); 
mux_module mux_module_inst_1_1199(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1201]),.i2(intermediate_reg_0[1200]),.o(intermediate_reg_1[600]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1200(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1199]),.i2(intermediate_reg_0[1198]),.o(intermediate_reg_1[599]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1201(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1197]),.i2(intermediate_reg_0[1196]),.o(intermediate_reg_1[598])); 
mux_module mux_module_inst_1_1202(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1195]),.i2(intermediate_reg_0[1194]),.o(intermediate_reg_1[597]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1203(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1193]),.i2(intermediate_reg_0[1192]),.o(intermediate_reg_1[596]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1204(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1191]),.i2(intermediate_reg_0[1190]),.o(intermediate_reg_1[595]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1205(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1189]),.i2(intermediate_reg_0[1188]),.o(intermediate_reg_1[594])); 
mux_module mux_module_inst_1_1206(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1187]),.i2(intermediate_reg_0[1186]),.o(intermediate_reg_1[593]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1207(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1185]),.i2(intermediate_reg_0[1184]),.o(intermediate_reg_1[592])); 
fsm fsm_inst_1_1208(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1183]),.i2(intermediate_reg_0[1182]),.o(intermediate_reg_1[591])); 
fsm fsm_inst_1_1209(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1181]),.i2(intermediate_reg_0[1180]),.o(intermediate_reg_1[590])); 
mux_module mux_module_inst_1_1210(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1179]),.i2(intermediate_reg_0[1178]),.o(intermediate_reg_1[589]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1211(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1177]),.i2(intermediate_reg_0[1176]),.o(intermediate_reg_1[588])); 
mux_module mux_module_inst_1_1212(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1175]),.i2(intermediate_reg_0[1174]),.o(intermediate_reg_1[587]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1213(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1173]),.i2(intermediate_reg_0[1172]),.o(intermediate_reg_1[586])); 
fsm fsm_inst_1_1214(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1171]),.i2(intermediate_reg_0[1170]),.o(intermediate_reg_1[585])); 
fsm fsm_inst_1_1215(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1169]),.i2(intermediate_reg_0[1168]),.o(intermediate_reg_1[584])); 
mux_module mux_module_inst_1_1216(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1167]),.i2(intermediate_reg_0[1166]),.o(intermediate_reg_1[583]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1217(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1165]),.i2(intermediate_reg_0[1164]),.o(intermediate_reg_1[582])); 
mux_module mux_module_inst_1_1218(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1163]),.i2(intermediate_reg_0[1162]),.o(intermediate_reg_1[581]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1219(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1161]),.i2(intermediate_reg_0[1160]),.o(intermediate_reg_1[580])); 
fsm fsm_inst_1_1220(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1159]),.i2(intermediate_reg_0[1158]),.o(intermediate_reg_1[579])); 
mux_module mux_module_inst_1_1221(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1157]),.i2(intermediate_reg_0[1156]),.o(intermediate_reg_1[578]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1222(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1155]),.i2(intermediate_reg_0[1154]),.o(intermediate_reg_1[577])); 
mux_module mux_module_inst_1_1223(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1153]),.i2(intermediate_reg_0[1152]),.o(intermediate_reg_1[576]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1224(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1151]),.i2(intermediate_reg_0[1150]),.o(intermediate_reg_1[575])); 
fsm fsm_inst_1_1225(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1149]),.i2(intermediate_reg_0[1148]),.o(intermediate_reg_1[574])); 
mux_module mux_module_inst_1_1226(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1147]),.i2(intermediate_reg_0[1146]),.o(intermediate_reg_1[573]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1227(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1145]),.i2(intermediate_reg_0[1144]),.o(intermediate_reg_1[572])); 
mux_module mux_module_inst_1_1228(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1143]),.i2(intermediate_reg_0[1142]),.o(intermediate_reg_1[571]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1229(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1141]),.i2(intermediate_reg_0[1140]),.o(intermediate_reg_1[570])); 
mux_module mux_module_inst_1_1230(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1139]),.i2(intermediate_reg_0[1138]),.o(intermediate_reg_1[569]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1231(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1137]),.i2(intermediate_reg_0[1136]),.o(intermediate_reg_1[568])); 
mux_module mux_module_inst_1_1232(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1135]),.i2(intermediate_reg_0[1134]),.o(intermediate_reg_1[567]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1233(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1133]),.i2(intermediate_reg_0[1132]),.o(intermediate_reg_1[566]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1234(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1131]),.i2(intermediate_reg_0[1130]),.o(intermediate_reg_1[565]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1235(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1129]),.i2(intermediate_reg_0[1128]),.o(intermediate_reg_1[564]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1236(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1127]),.i2(intermediate_reg_0[1126]),.o(intermediate_reg_1[563]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1237(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1125]),.i2(intermediate_reg_0[1124]),.o(intermediate_reg_1[562])); 
fsm fsm_inst_1_1238(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1123]),.i2(intermediate_reg_0[1122]),.o(intermediate_reg_1[561])); 
mux_module mux_module_inst_1_1239(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1121]),.i2(intermediate_reg_0[1120]),.o(intermediate_reg_1[560]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1240(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1119]),.i2(intermediate_reg_0[1118]),.o(intermediate_reg_1[559]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1241(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1117]),.i2(intermediate_reg_0[1116]),.o(intermediate_reg_1[558])); 
fsm fsm_inst_1_1242(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1115]),.i2(intermediate_reg_0[1114]),.o(intermediate_reg_1[557])); 
fsm fsm_inst_1_1243(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1113]),.i2(intermediate_reg_0[1112]),.o(intermediate_reg_1[556])); 
fsm fsm_inst_1_1244(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1111]),.i2(intermediate_reg_0[1110]),.o(intermediate_reg_1[555])); 
fsm fsm_inst_1_1245(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1109]),.i2(intermediate_reg_0[1108]),.o(intermediate_reg_1[554])); 
fsm fsm_inst_1_1246(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1107]),.i2(intermediate_reg_0[1106]),.o(intermediate_reg_1[553])); 
fsm fsm_inst_1_1247(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1105]),.i2(intermediate_reg_0[1104]),.o(intermediate_reg_1[552])); 
mux_module mux_module_inst_1_1248(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1103]),.i2(intermediate_reg_0[1102]),.o(intermediate_reg_1[551]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1249(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1101]),.i2(intermediate_reg_0[1100]),.o(intermediate_reg_1[550]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1250(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1099]),.i2(intermediate_reg_0[1098]),.o(intermediate_reg_1[549]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1251(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1097]),.i2(intermediate_reg_0[1096]),.o(intermediate_reg_1[548]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1252(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1095]),.i2(intermediate_reg_0[1094]),.o(intermediate_reg_1[547]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1253(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1093]),.i2(intermediate_reg_0[1092]),.o(intermediate_reg_1[546]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1254(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1091]),.i2(intermediate_reg_0[1090]),.o(intermediate_reg_1[545]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1255(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1089]),.i2(intermediate_reg_0[1088]),.o(intermediate_reg_1[544])); 
fsm fsm_inst_1_1256(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1087]),.i2(intermediate_reg_0[1086]),.o(intermediate_reg_1[543])); 
mux_module mux_module_inst_1_1257(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1085]),.i2(intermediate_reg_0[1084]),.o(intermediate_reg_1[542]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1258(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1083]),.i2(intermediate_reg_0[1082]),.o(intermediate_reg_1[541])); 
fsm fsm_inst_1_1259(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1081]),.i2(intermediate_reg_0[1080]),.o(intermediate_reg_1[540])); 
mux_module mux_module_inst_1_1260(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1079]),.i2(intermediate_reg_0[1078]),.o(intermediate_reg_1[539]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1261(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1077]),.i2(intermediate_reg_0[1076]),.o(intermediate_reg_1[538]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1262(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1075]),.i2(intermediate_reg_0[1074]),.o(intermediate_reg_1[537]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1263(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1073]),.i2(intermediate_reg_0[1072]),.o(intermediate_reg_1[536]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1264(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1071]),.i2(intermediate_reg_0[1070]),.o(intermediate_reg_1[535]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1265(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1069]),.i2(intermediate_reg_0[1068]),.o(intermediate_reg_1[534]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1266(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1067]),.i2(intermediate_reg_0[1066]),.o(intermediate_reg_1[533])); 
mux_module mux_module_inst_1_1267(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1065]),.i2(intermediate_reg_0[1064]),.o(intermediate_reg_1[532]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1268(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1063]),.i2(intermediate_reg_0[1062]),.o(intermediate_reg_1[531]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1269(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1061]),.i2(intermediate_reg_0[1060]),.o(intermediate_reg_1[530]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1270(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1059]),.i2(intermediate_reg_0[1058]),.o(intermediate_reg_1[529]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1271(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1057]),.i2(intermediate_reg_0[1056]),.o(intermediate_reg_1[528]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1272(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1055]),.i2(intermediate_reg_0[1054]),.o(intermediate_reg_1[527]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1273(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1053]),.i2(intermediate_reg_0[1052]),.o(intermediate_reg_1[526])); 
fsm fsm_inst_1_1274(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1051]),.i2(intermediate_reg_0[1050]),.o(intermediate_reg_1[525])); 
mux_module mux_module_inst_1_1275(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1049]),.i2(intermediate_reg_0[1048]),.o(intermediate_reg_1[524]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1276(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1047]),.i2(intermediate_reg_0[1046]),.o(intermediate_reg_1[523]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1277(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1045]),.i2(intermediate_reg_0[1044]),.o(intermediate_reg_1[522]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1278(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1043]),.i2(intermediate_reg_0[1042]),.o(intermediate_reg_1[521])); 
mux_module mux_module_inst_1_1279(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1041]),.i2(intermediate_reg_0[1040]),.o(intermediate_reg_1[520]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1280(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1039]),.i2(intermediate_reg_0[1038]),.o(intermediate_reg_1[519]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1281(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1037]),.i2(intermediate_reg_0[1036]),.o(intermediate_reg_1[518])); 
fsm fsm_inst_1_1282(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1035]),.i2(intermediate_reg_0[1034]),.o(intermediate_reg_1[517])); 
mux_module mux_module_inst_1_1283(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1033]),.i2(intermediate_reg_0[1032]),.o(intermediate_reg_1[516]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1284(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1031]),.i2(intermediate_reg_0[1030]),.o(intermediate_reg_1[515])); 
fsm fsm_inst_1_1285(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1029]),.i2(intermediate_reg_0[1028]),.o(intermediate_reg_1[514])); 
mux_module mux_module_inst_1_1286(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1027]),.i2(intermediate_reg_0[1026]),.o(intermediate_reg_1[513]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1287(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1025]),.i2(intermediate_reg_0[1024]),.o(intermediate_reg_1[512])); 
fsm fsm_inst_1_1288(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1023]),.i2(intermediate_reg_0[1022]),.o(intermediate_reg_1[511])); 
mux_module mux_module_inst_1_1289(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1021]),.i2(intermediate_reg_0[1020]),.o(intermediate_reg_1[510]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1290(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1019]),.i2(intermediate_reg_0[1018]),.o(intermediate_reg_1[509]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1291(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1017]),.i2(intermediate_reg_0[1016]),.o(intermediate_reg_1[508]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1292(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1015]),.i2(intermediate_reg_0[1014]),.o(intermediate_reg_1[507])); 
mux_module mux_module_inst_1_1293(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1013]),.i2(intermediate_reg_0[1012]),.o(intermediate_reg_1[506]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1294(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1011]),.i2(intermediate_reg_0[1010]),.o(intermediate_reg_1[505])); 
mux_module mux_module_inst_1_1295(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1009]),.i2(intermediate_reg_0[1008]),.o(intermediate_reg_1[504]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1296(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1007]),.i2(intermediate_reg_0[1006]),.o(intermediate_reg_1[503]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1297(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1005]),.i2(intermediate_reg_0[1004]),.o(intermediate_reg_1[502]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1298(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1003]),.i2(intermediate_reg_0[1002]),.o(intermediate_reg_1[501]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1299(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1001]),.i2(intermediate_reg_0[1000]),.o(intermediate_reg_1[500])); 
mux_module mux_module_inst_1_1300(.clk(clk),.reset(reset),.i1(intermediate_reg_0[999]),.i2(intermediate_reg_0[998]),.o(intermediate_reg_1[499]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1301(.clk(clk),.reset(reset),.i1(intermediate_reg_0[997]),.i2(intermediate_reg_0[996]),.o(intermediate_reg_1[498])); 
mux_module mux_module_inst_1_1302(.clk(clk),.reset(reset),.i1(intermediate_reg_0[995]),.i2(intermediate_reg_0[994]),.o(intermediate_reg_1[497]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1303(.clk(clk),.reset(reset),.i1(intermediate_reg_0[993]),.i2(intermediate_reg_0[992]),.o(intermediate_reg_1[496])); 
fsm fsm_inst_1_1304(.clk(clk),.reset(reset),.i1(intermediate_reg_0[991]),.i2(intermediate_reg_0[990]),.o(intermediate_reg_1[495])); 
fsm fsm_inst_1_1305(.clk(clk),.reset(reset),.i1(intermediate_reg_0[989]),.i2(intermediate_reg_0[988]),.o(intermediate_reg_1[494])); 
mux_module mux_module_inst_1_1306(.clk(clk),.reset(reset),.i1(intermediate_reg_0[987]),.i2(intermediate_reg_0[986]),.o(intermediate_reg_1[493]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1307(.clk(clk),.reset(reset),.i1(intermediate_reg_0[985]),.i2(intermediate_reg_0[984]),.o(intermediate_reg_1[492]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1308(.clk(clk),.reset(reset),.i1(intermediate_reg_0[983]),.i2(intermediate_reg_0[982]),.o(intermediate_reg_1[491]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1309(.clk(clk),.reset(reset),.i1(intermediate_reg_0[981]),.i2(intermediate_reg_0[980]),.o(intermediate_reg_1[490]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1310(.clk(clk),.reset(reset),.i1(intermediate_reg_0[979]),.i2(intermediate_reg_0[978]),.o(intermediate_reg_1[489])); 
mux_module mux_module_inst_1_1311(.clk(clk),.reset(reset),.i1(intermediate_reg_0[977]),.i2(intermediate_reg_0[976]),.o(intermediate_reg_1[488]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1312(.clk(clk),.reset(reset),.i1(intermediate_reg_0[975]),.i2(intermediate_reg_0[974]),.o(intermediate_reg_1[487]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1313(.clk(clk),.reset(reset),.i1(intermediate_reg_0[973]),.i2(intermediate_reg_0[972]),.o(intermediate_reg_1[486]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1314(.clk(clk),.reset(reset),.i1(intermediate_reg_0[971]),.i2(intermediate_reg_0[970]),.o(intermediate_reg_1[485])); 
fsm fsm_inst_1_1315(.clk(clk),.reset(reset),.i1(intermediate_reg_0[969]),.i2(intermediate_reg_0[968]),.o(intermediate_reg_1[484])); 
fsm fsm_inst_1_1316(.clk(clk),.reset(reset),.i1(intermediate_reg_0[967]),.i2(intermediate_reg_0[966]),.o(intermediate_reg_1[483])); 
mux_module mux_module_inst_1_1317(.clk(clk),.reset(reset),.i1(intermediate_reg_0[965]),.i2(intermediate_reg_0[964]),.o(intermediate_reg_1[482]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1318(.clk(clk),.reset(reset),.i1(intermediate_reg_0[963]),.i2(intermediate_reg_0[962]),.o(intermediate_reg_1[481])); 
fsm fsm_inst_1_1319(.clk(clk),.reset(reset),.i1(intermediate_reg_0[961]),.i2(intermediate_reg_0[960]),.o(intermediate_reg_1[480])); 
fsm fsm_inst_1_1320(.clk(clk),.reset(reset),.i1(intermediate_reg_0[959]),.i2(intermediate_reg_0[958]),.o(intermediate_reg_1[479])); 
fsm fsm_inst_1_1321(.clk(clk),.reset(reset),.i1(intermediate_reg_0[957]),.i2(intermediate_reg_0[956]),.o(intermediate_reg_1[478])); 
fsm fsm_inst_1_1322(.clk(clk),.reset(reset),.i1(intermediate_reg_0[955]),.i2(intermediate_reg_0[954]),.o(intermediate_reg_1[477])); 
fsm fsm_inst_1_1323(.clk(clk),.reset(reset),.i1(intermediate_reg_0[953]),.i2(intermediate_reg_0[952]),.o(intermediate_reg_1[476])); 
mux_module mux_module_inst_1_1324(.clk(clk),.reset(reset),.i1(intermediate_reg_0[951]),.i2(intermediate_reg_0[950]),.o(intermediate_reg_1[475]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1325(.clk(clk),.reset(reset),.i1(intermediate_reg_0[949]),.i2(intermediate_reg_0[948]),.o(intermediate_reg_1[474]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1326(.clk(clk),.reset(reset),.i1(intermediate_reg_0[947]),.i2(intermediate_reg_0[946]),.o(intermediate_reg_1[473])); 
fsm fsm_inst_1_1327(.clk(clk),.reset(reset),.i1(intermediate_reg_0[945]),.i2(intermediate_reg_0[944]),.o(intermediate_reg_1[472])); 
mux_module mux_module_inst_1_1328(.clk(clk),.reset(reset),.i1(intermediate_reg_0[943]),.i2(intermediate_reg_0[942]),.o(intermediate_reg_1[471]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1329(.clk(clk),.reset(reset),.i1(intermediate_reg_0[941]),.i2(intermediate_reg_0[940]),.o(intermediate_reg_1[470])); 
mux_module mux_module_inst_1_1330(.clk(clk),.reset(reset),.i1(intermediate_reg_0[939]),.i2(intermediate_reg_0[938]),.o(intermediate_reg_1[469]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1331(.clk(clk),.reset(reset),.i1(intermediate_reg_0[937]),.i2(intermediate_reg_0[936]),.o(intermediate_reg_1[468]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1332(.clk(clk),.reset(reset),.i1(intermediate_reg_0[935]),.i2(intermediate_reg_0[934]),.o(intermediate_reg_1[467])); 
fsm fsm_inst_1_1333(.clk(clk),.reset(reset),.i1(intermediate_reg_0[933]),.i2(intermediate_reg_0[932]),.o(intermediate_reg_1[466])); 
fsm fsm_inst_1_1334(.clk(clk),.reset(reset),.i1(intermediate_reg_0[931]),.i2(intermediate_reg_0[930]),.o(intermediate_reg_1[465])); 
fsm fsm_inst_1_1335(.clk(clk),.reset(reset),.i1(intermediate_reg_0[929]),.i2(intermediate_reg_0[928]),.o(intermediate_reg_1[464])); 
fsm fsm_inst_1_1336(.clk(clk),.reset(reset),.i1(intermediate_reg_0[927]),.i2(intermediate_reg_0[926]),.o(intermediate_reg_1[463])); 
mux_module mux_module_inst_1_1337(.clk(clk),.reset(reset),.i1(intermediate_reg_0[925]),.i2(intermediate_reg_0[924]),.o(intermediate_reg_1[462]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1338(.clk(clk),.reset(reset),.i1(intermediate_reg_0[923]),.i2(intermediate_reg_0[922]),.o(intermediate_reg_1[461]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1339(.clk(clk),.reset(reset),.i1(intermediate_reg_0[921]),.i2(intermediate_reg_0[920]),.o(intermediate_reg_1[460]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1340(.clk(clk),.reset(reset),.i1(intermediate_reg_0[919]),.i2(intermediate_reg_0[918]),.o(intermediate_reg_1[459])); 
mux_module mux_module_inst_1_1341(.clk(clk),.reset(reset),.i1(intermediate_reg_0[917]),.i2(intermediate_reg_0[916]),.o(intermediate_reg_1[458]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1342(.clk(clk),.reset(reset),.i1(intermediate_reg_0[915]),.i2(intermediate_reg_0[914]),.o(intermediate_reg_1[457]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1343(.clk(clk),.reset(reset),.i1(intermediate_reg_0[913]),.i2(intermediate_reg_0[912]),.o(intermediate_reg_1[456])); 
fsm fsm_inst_1_1344(.clk(clk),.reset(reset),.i1(intermediate_reg_0[911]),.i2(intermediate_reg_0[910]),.o(intermediate_reg_1[455])); 
fsm fsm_inst_1_1345(.clk(clk),.reset(reset),.i1(intermediate_reg_0[909]),.i2(intermediate_reg_0[908]),.o(intermediate_reg_1[454])); 
mux_module mux_module_inst_1_1346(.clk(clk),.reset(reset),.i1(intermediate_reg_0[907]),.i2(intermediate_reg_0[906]),.o(intermediate_reg_1[453]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1347(.clk(clk),.reset(reset),.i1(intermediate_reg_0[905]),.i2(intermediate_reg_0[904]),.o(intermediate_reg_1[452])); 
mux_module mux_module_inst_1_1348(.clk(clk),.reset(reset),.i1(intermediate_reg_0[903]),.i2(intermediate_reg_0[902]),.o(intermediate_reg_1[451]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1349(.clk(clk),.reset(reset),.i1(intermediate_reg_0[901]),.i2(intermediate_reg_0[900]),.o(intermediate_reg_1[450]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1350(.clk(clk),.reset(reset),.i1(intermediate_reg_0[899]),.i2(intermediate_reg_0[898]),.o(intermediate_reg_1[449]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1351(.clk(clk),.reset(reset),.i1(intermediate_reg_0[897]),.i2(intermediate_reg_0[896]),.o(intermediate_reg_1[448]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1352(.clk(clk),.reset(reset),.i1(intermediate_reg_0[895]),.i2(intermediate_reg_0[894]),.o(intermediate_reg_1[447]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1353(.clk(clk),.reset(reset),.i1(intermediate_reg_0[893]),.i2(intermediate_reg_0[892]),.o(intermediate_reg_1[446])); 
fsm fsm_inst_1_1354(.clk(clk),.reset(reset),.i1(intermediate_reg_0[891]),.i2(intermediate_reg_0[890]),.o(intermediate_reg_1[445])); 
fsm fsm_inst_1_1355(.clk(clk),.reset(reset),.i1(intermediate_reg_0[889]),.i2(intermediate_reg_0[888]),.o(intermediate_reg_1[444])); 
fsm fsm_inst_1_1356(.clk(clk),.reset(reset),.i1(intermediate_reg_0[887]),.i2(intermediate_reg_0[886]),.o(intermediate_reg_1[443])); 
fsm fsm_inst_1_1357(.clk(clk),.reset(reset),.i1(intermediate_reg_0[885]),.i2(intermediate_reg_0[884]),.o(intermediate_reg_1[442])); 
fsm fsm_inst_1_1358(.clk(clk),.reset(reset),.i1(intermediate_reg_0[883]),.i2(intermediate_reg_0[882]),.o(intermediate_reg_1[441])); 
mux_module mux_module_inst_1_1359(.clk(clk),.reset(reset),.i1(intermediate_reg_0[881]),.i2(intermediate_reg_0[880]),.o(intermediate_reg_1[440]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1360(.clk(clk),.reset(reset),.i1(intermediate_reg_0[879]),.i2(intermediate_reg_0[878]),.o(intermediate_reg_1[439])); 
fsm fsm_inst_1_1361(.clk(clk),.reset(reset),.i1(intermediate_reg_0[877]),.i2(intermediate_reg_0[876]),.o(intermediate_reg_1[438])); 
mux_module mux_module_inst_1_1362(.clk(clk),.reset(reset),.i1(intermediate_reg_0[875]),.i2(intermediate_reg_0[874]),.o(intermediate_reg_1[437]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1363(.clk(clk),.reset(reset),.i1(intermediate_reg_0[873]),.i2(intermediate_reg_0[872]),.o(intermediate_reg_1[436]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1364(.clk(clk),.reset(reset),.i1(intermediate_reg_0[871]),.i2(intermediate_reg_0[870]),.o(intermediate_reg_1[435])); 
fsm fsm_inst_1_1365(.clk(clk),.reset(reset),.i1(intermediate_reg_0[869]),.i2(intermediate_reg_0[868]),.o(intermediate_reg_1[434])); 
mux_module mux_module_inst_1_1366(.clk(clk),.reset(reset),.i1(intermediate_reg_0[867]),.i2(intermediate_reg_0[866]),.o(intermediate_reg_1[433]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1367(.clk(clk),.reset(reset),.i1(intermediate_reg_0[865]),.i2(intermediate_reg_0[864]),.o(intermediate_reg_1[432])); 
fsm fsm_inst_1_1368(.clk(clk),.reset(reset),.i1(intermediate_reg_0[863]),.i2(intermediate_reg_0[862]),.o(intermediate_reg_1[431])); 
mux_module mux_module_inst_1_1369(.clk(clk),.reset(reset),.i1(intermediate_reg_0[861]),.i2(intermediate_reg_0[860]),.o(intermediate_reg_1[430]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1370(.clk(clk),.reset(reset),.i1(intermediate_reg_0[859]),.i2(intermediate_reg_0[858]),.o(intermediate_reg_1[429])); 
fsm fsm_inst_1_1371(.clk(clk),.reset(reset),.i1(intermediate_reg_0[857]),.i2(intermediate_reg_0[856]),.o(intermediate_reg_1[428])); 
fsm fsm_inst_1_1372(.clk(clk),.reset(reset),.i1(intermediate_reg_0[855]),.i2(intermediate_reg_0[854]),.o(intermediate_reg_1[427])); 
fsm fsm_inst_1_1373(.clk(clk),.reset(reset),.i1(intermediate_reg_0[853]),.i2(intermediate_reg_0[852]),.o(intermediate_reg_1[426])); 
mux_module mux_module_inst_1_1374(.clk(clk),.reset(reset),.i1(intermediate_reg_0[851]),.i2(intermediate_reg_0[850]),.o(intermediate_reg_1[425]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1375(.clk(clk),.reset(reset),.i1(intermediate_reg_0[849]),.i2(intermediate_reg_0[848]),.o(intermediate_reg_1[424]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1376(.clk(clk),.reset(reset),.i1(intermediate_reg_0[847]),.i2(intermediate_reg_0[846]),.o(intermediate_reg_1[423])); 
fsm fsm_inst_1_1377(.clk(clk),.reset(reset),.i1(intermediate_reg_0[845]),.i2(intermediate_reg_0[844]),.o(intermediate_reg_1[422])); 
fsm fsm_inst_1_1378(.clk(clk),.reset(reset),.i1(intermediate_reg_0[843]),.i2(intermediate_reg_0[842]),.o(intermediate_reg_1[421])); 
mux_module mux_module_inst_1_1379(.clk(clk),.reset(reset),.i1(intermediate_reg_0[841]),.i2(intermediate_reg_0[840]),.o(intermediate_reg_1[420]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1380(.clk(clk),.reset(reset),.i1(intermediate_reg_0[839]),.i2(intermediate_reg_0[838]),.o(intermediate_reg_1[419]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1381(.clk(clk),.reset(reset),.i1(intermediate_reg_0[837]),.i2(intermediate_reg_0[836]),.o(intermediate_reg_1[418]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1382(.clk(clk),.reset(reset),.i1(intermediate_reg_0[835]),.i2(intermediate_reg_0[834]),.o(intermediate_reg_1[417])); 
fsm fsm_inst_1_1383(.clk(clk),.reset(reset),.i1(intermediate_reg_0[833]),.i2(intermediate_reg_0[832]),.o(intermediate_reg_1[416])); 
fsm fsm_inst_1_1384(.clk(clk),.reset(reset),.i1(intermediate_reg_0[831]),.i2(intermediate_reg_0[830]),.o(intermediate_reg_1[415])); 
mux_module mux_module_inst_1_1385(.clk(clk),.reset(reset),.i1(intermediate_reg_0[829]),.i2(intermediate_reg_0[828]),.o(intermediate_reg_1[414]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1386(.clk(clk),.reset(reset),.i1(intermediate_reg_0[827]),.i2(intermediate_reg_0[826]),.o(intermediate_reg_1[413]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1387(.clk(clk),.reset(reset),.i1(intermediate_reg_0[825]),.i2(intermediate_reg_0[824]),.o(intermediate_reg_1[412])); 
fsm fsm_inst_1_1388(.clk(clk),.reset(reset),.i1(intermediate_reg_0[823]),.i2(intermediate_reg_0[822]),.o(intermediate_reg_1[411])); 
fsm fsm_inst_1_1389(.clk(clk),.reset(reset),.i1(intermediate_reg_0[821]),.i2(intermediate_reg_0[820]),.o(intermediate_reg_1[410])); 
mux_module mux_module_inst_1_1390(.clk(clk),.reset(reset),.i1(intermediate_reg_0[819]),.i2(intermediate_reg_0[818]),.o(intermediate_reg_1[409]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1391(.clk(clk),.reset(reset),.i1(intermediate_reg_0[817]),.i2(intermediate_reg_0[816]),.o(intermediate_reg_1[408])); 
mux_module mux_module_inst_1_1392(.clk(clk),.reset(reset),.i1(intermediate_reg_0[815]),.i2(intermediate_reg_0[814]),.o(intermediate_reg_1[407]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1393(.clk(clk),.reset(reset),.i1(intermediate_reg_0[813]),.i2(intermediate_reg_0[812]),.o(intermediate_reg_1[406])); 
mux_module mux_module_inst_1_1394(.clk(clk),.reset(reset),.i1(intermediate_reg_0[811]),.i2(intermediate_reg_0[810]),.o(intermediate_reg_1[405]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1395(.clk(clk),.reset(reset),.i1(intermediate_reg_0[809]),.i2(intermediate_reg_0[808]),.o(intermediate_reg_1[404]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1396(.clk(clk),.reset(reset),.i1(intermediate_reg_0[807]),.i2(intermediate_reg_0[806]),.o(intermediate_reg_1[403])); 
mux_module mux_module_inst_1_1397(.clk(clk),.reset(reset),.i1(intermediate_reg_0[805]),.i2(intermediate_reg_0[804]),.o(intermediate_reg_1[402]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1398(.clk(clk),.reset(reset),.i1(intermediate_reg_0[803]),.i2(intermediate_reg_0[802]),.o(intermediate_reg_1[401]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1399(.clk(clk),.reset(reset),.i1(intermediate_reg_0[801]),.i2(intermediate_reg_0[800]),.o(intermediate_reg_1[400])); 
fsm fsm_inst_1_1400(.clk(clk),.reset(reset),.i1(intermediate_reg_0[799]),.i2(intermediate_reg_0[798]),.o(intermediate_reg_1[399])); 
fsm fsm_inst_1_1401(.clk(clk),.reset(reset),.i1(intermediate_reg_0[797]),.i2(intermediate_reg_0[796]),.o(intermediate_reg_1[398])); 
fsm fsm_inst_1_1402(.clk(clk),.reset(reset),.i1(intermediate_reg_0[795]),.i2(intermediate_reg_0[794]),.o(intermediate_reg_1[397])); 
fsm fsm_inst_1_1403(.clk(clk),.reset(reset),.i1(intermediate_reg_0[793]),.i2(intermediate_reg_0[792]),.o(intermediate_reg_1[396])); 
mux_module mux_module_inst_1_1404(.clk(clk),.reset(reset),.i1(intermediate_reg_0[791]),.i2(intermediate_reg_0[790]),.o(intermediate_reg_1[395]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1405(.clk(clk),.reset(reset),.i1(intermediate_reg_0[789]),.i2(intermediate_reg_0[788]),.o(intermediate_reg_1[394])); 
fsm fsm_inst_1_1406(.clk(clk),.reset(reset),.i1(intermediate_reg_0[787]),.i2(intermediate_reg_0[786]),.o(intermediate_reg_1[393])); 
mux_module mux_module_inst_1_1407(.clk(clk),.reset(reset),.i1(intermediate_reg_0[785]),.i2(intermediate_reg_0[784]),.o(intermediate_reg_1[392]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1408(.clk(clk),.reset(reset),.i1(intermediate_reg_0[783]),.i2(intermediate_reg_0[782]),.o(intermediate_reg_1[391])); 
mux_module mux_module_inst_1_1409(.clk(clk),.reset(reset),.i1(intermediate_reg_0[781]),.i2(intermediate_reg_0[780]),.o(intermediate_reg_1[390]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1410(.clk(clk),.reset(reset),.i1(intermediate_reg_0[779]),.i2(intermediate_reg_0[778]),.o(intermediate_reg_1[389])); 
fsm fsm_inst_1_1411(.clk(clk),.reset(reset),.i1(intermediate_reg_0[777]),.i2(intermediate_reg_0[776]),.o(intermediate_reg_1[388])); 
mux_module mux_module_inst_1_1412(.clk(clk),.reset(reset),.i1(intermediate_reg_0[775]),.i2(intermediate_reg_0[774]),.o(intermediate_reg_1[387]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1413(.clk(clk),.reset(reset),.i1(intermediate_reg_0[773]),.i2(intermediate_reg_0[772]),.o(intermediate_reg_1[386]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1414(.clk(clk),.reset(reset),.i1(intermediate_reg_0[771]),.i2(intermediate_reg_0[770]),.o(intermediate_reg_1[385])); 
mux_module mux_module_inst_1_1415(.clk(clk),.reset(reset),.i1(intermediate_reg_0[769]),.i2(intermediate_reg_0[768]),.o(intermediate_reg_1[384]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1416(.clk(clk),.reset(reset),.i1(intermediate_reg_0[767]),.i2(intermediate_reg_0[766]),.o(intermediate_reg_1[383])); 
mux_module mux_module_inst_1_1417(.clk(clk),.reset(reset),.i1(intermediate_reg_0[765]),.i2(intermediate_reg_0[764]),.o(intermediate_reg_1[382]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1418(.clk(clk),.reset(reset),.i1(intermediate_reg_0[763]),.i2(intermediate_reg_0[762]),.o(intermediate_reg_1[381])); 
mux_module mux_module_inst_1_1419(.clk(clk),.reset(reset),.i1(intermediate_reg_0[761]),.i2(intermediate_reg_0[760]),.o(intermediate_reg_1[380]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1420(.clk(clk),.reset(reset),.i1(intermediate_reg_0[759]),.i2(intermediate_reg_0[758]),.o(intermediate_reg_1[379])); 
fsm fsm_inst_1_1421(.clk(clk),.reset(reset),.i1(intermediate_reg_0[757]),.i2(intermediate_reg_0[756]),.o(intermediate_reg_1[378])); 
fsm fsm_inst_1_1422(.clk(clk),.reset(reset),.i1(intermediate_reg_0[755]),.i2(intermediate_reg_0[754]),.o(intermediate_reg_1[377])); 
fsm fsm_inst_1_1423(.clk(clk),.reset(reset),.i1(intermediate_reg_0[753]),.i2(intermediate_reg_0[752]),.o(intermediate_reg_1[376])); 
mux_module mux_module_inst_1_1424(.clk(clk),.reset(reset),.i1(intermediate_reg_0[751]),.i2(intermediate_reg_0[750]),.o(intermediate_reg_1[375]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1425(.clk(clk),.reset(reset),.i1(intermediate_reg_0[749]),.i2(intermediate_reg_0[748]),.o(intermediate_reg_1[374])); 
mux_module mux_module_inst_1_1426(.clk(clk),.reset(reset),.i1(intermediate_reg_0[747]),.i2(intermediate_reg_0[746]),.o(intermediate_reg_1[373]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1427(.clk(clk),.reset(reset),.i1(intermediate_reg_0[745]),.i2(intermediate_reg_0[744]),.o(intermediate_reg_1[372])); 
mux_module mux_module_inst_1_1428(.clk(clk),.reset(reset),.i1(intermediate_reg_0[743]),.i2(intermediate_reg_0[742]),.o(intermediate_reg_1[371]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1429(.clk(clk),.reset(reset),.i1(intermediate_reg_0[741]),.i2(intermediate_reg_0[740]),.o(intermediate_reg_1[370]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1430(.clk(clk),.reset(reset),.i1(intermediate_reg_0[739]),.i2(intermediate_reg_0[738]),.o(intermediate_reg_1[369])); 
mux_module mux_module_inst_1_1431(.clk(clk),.reset(reset),.i1(intermediate_reg_0[737]),.i2(intermediate_reg_0[736]),.o(intermediate_reg_1[368]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1432(.clk(clk),.reset(reset),.i1(intermediate_reg_0[735]),.i2(intermediate_reg_0[734]),.o(intermediate_reg_1[367])); 
fsm fsm_inst_1_1433(.clk(clk),.reset(reset),.i1(intermediate_reg_0[733]),.i2(intermediate_reg_0[732]),.o(intermediate_reg_1[366])); 
mux_module mux_module_inst_1_1434(.clk(clk),.reset(reset),.i1(intermediate_reg_0[731]),.i2(intermediate_reg_0[730]),.o(intermediate_reg_1[365]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1435(.clk(clk),.reset(reset),.i1(intermediate_reg_0[729]),.i2(intermediate_reg_0[728]),.o(intermediate_reg_1[364]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1436(.clk(clk),.reset(reset),.i1(intermediate_reg_0[727]),.i2(intermediate_reg_0[726]),.o(intermediate_reg_1[363])); 
fsm fsm_inst_1_1437(.clk(clk),.reset(reset),.i1(intermediate_reg_0[725]),.i2(intermediate_reg_0[724]),.o(intermediate_reg_1[362])); 
mux_module mux_module_inst_1_1438(.clk(clk),.reset(reset),.i1(intermediate_reg_0[723]),.i2(intermediate_reg_0[722]),.o(intermediate_reg_1[361]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1439(.clk(clk),.reset(reset),.i1(intermediate_reg_0[721]),.i2(intermediate_reg_0[720]),.o(intermediate_reg_1[360]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1440(.clk(clk),.reset(reset),.i1(intermediate_reg_0[719]),.i2(intermediate_reg_0[718]),.o(intermediate_reg_1[359]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1441(.clk(clk),.reset(reset),.i1(intermediate_reg_0[717]),.i2(intermediate_reg_0[716]),.o(intermediate_reg_1[358]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1442(.clk(clk),.reset(reset),.i1(intermediate_reg_0[715]),.i2(intermediate_reg_0[714]),.o(intermediate_reg_1[357]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1443(.clk(clk),.reset(reset),.i1(intermediate_reg_0[713]),.i2(intermediate_reg_0[712]),.o(intermediate_reg_1[356])); 
fsm fsm_inst_1_1444(.clk(clk),.reset(reset),.i1(intermediate_reg_0[711]),.i2(intermediate_reg_0[710]),.o(intermediate_reg_1[355])); 
mux_module mux_module_inst_1_1445(.clk(clk),.reset(reset),.i1(intermediate_reg_0[709]),.i2(intermediate_reg_0[708]),.o(intermediate_reg_1[354]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1446(.clk(clk),.reset(reset),.i1(intermediate_reg_0[707]),.i2(intermediate_reg_0[706]),.o(intermediate_reg_1[353])); 
mux_module mux_module_inst_1_1447(.clk(clk),.reset(reset),.i1(intermediate_reg_0[705]),.i2(intermediate_reg_0[704]),.o(intermediate_reg_1[352]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1448(.clk(clk),.reset(reset),.i1(intermediate_reg_0[703]),.i2(intermediate_reg_0[702]),.o(intermediate_reg_1[351]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1449(.clk(clk),.reset(reset),.i1(intermediate_reg_0[701]),.i2(intermediate_reg_0[700]),.o(intermediate_reg_1[350]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1450(.clk(clk),.reset(reset),.i1(intermediate_reg_0[699]),.i2(intermediate_reg_0[698]),.o(intermediate_reg_1[349]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1451(.clk(clk),.reset(reset),.i1(intermediate_reg_0[697]),.i2(intermediate_reg_0[696]),.o(intermediate_reg_1[348])); 
mux_module mux_module_inst_1_1452(.clk(clk),.reset(reset),.i1(intermediate_reg_0[695]),.i2(intermediate_reg_0[694]),.o(intermediate_reg_1[347]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1453(.clk(clk),.reset(reset),.i1(intermediate_reg_0[693]),.i2(intermediate_reg_0[692]),.o(intermediate_reg_1[346]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1454(.clk(clk),.reset(reset),.i1(intermediate_reg_0[691]),.i2(intermediate_reg_0[690]),.o(intermediate_reg_1[345]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1455(.clk(clk),.reset(reset),.i1(intermediate_reg_0[689]),.i2(intermediate_reg_0[688]),.o(intermediate_reg_1[344]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1456(.clk(clk),.reset(reset),.i1(intermediate_reg_0[687]),.i2(intermediate_reg_0[686]),.o(intermediate_reg_1[343])); 
mux_module mux_module_inst_1_1457(.clk(clk),.reset(reset),.i1(intermediate_reg_0[685]),.i2(intermediate_reg_0[684]),.o(intermediate_reg_1[342]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1458(.clk(clk),.reset(reset),.i1(intermediate_reg_0[683]),.i2(intermediate_reg_0[682]),.o(intermediate_reg_1[341]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1459(.clk(clk),.reset(reset),.i1(intermediate_reg_0[681]),.i2(intermediate_reg_0[680]),.o(intermediate_reg_1[340])); 
mux_module mux_module_inst_1_1460(.clk(clk),.reset(reset),.i1(intermediate_reg_0[679]),.i2(intermediate_reg_0[678]),.o(intermediate_reg_1[339]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1461(.clk(clk),.reset(reset),.i1(intermediate_reg_0[677]),.i2(intermediate_reg_0[676]),.o(intermediate_reg_1[338]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1462(.clk(clk),.reset(reset),.i1(intermediate_reg_0[675]),.i2(intermediate_reg_0[674]),.o(intermediate_reg_1[337]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1463(.clk(clk),.reset(reset),.i1(intermediate_reg_0[673]),.i2(intermediate_reg_0[672]),.o(intermediate_reg_1[336])); 
mux_module mux_module_inst_1_1464(.clk(clk),.reset(reset),.i1(intermediate_reg_0[671]),.i2(intermediate_reg_0[670]),.o(intermediate_reg_1[335]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1465(.clk(clk),.reset(reset),.i1(intermediate_reg_0[669]),.i2(intermediate_reg_0[668]),.o(intermediate_reg_1[334])); 
fsm fsm_inst_1_1466(.clk(clk),.reset(reset),.i1(intermediate_reg_0[667]),.i2(intermediate_reg_0[666]),.o(intermediate_reg_1[333])); 
fsm fsm_inst_1_1467(.clk(clk),.reset(reset),.i1(intermediate_reg_0[665]),.i2(intermediate_reg_0[664]),.o(intermediate_reg_1[332])); 
fsm fsm_inst_1_1468(.clk(clk),.reset(reset),.i1(intermediate_reg_0[663]),.i2(intermediate_reg_0[662]),.o(intermediate_reg_1[331])); 
mux_module mux_module_inst_1_1469(.clk(clk),.reset(reset),.i1(intermediate_reg_0[661]),.i2(intermediate_reg_0[660]),.o(intermediate_reg_1[330]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1470(.clk(clk),.reset(reset),.i1(intermediate_reg_0[659]),.i2(intermediate_reg_0[658]),.o(intermediate_reg_1[329]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1471(.clk(clk),.reset(reset),.i1(intermediate_reg_0[657]),.i2(intermediate_reg_0[656]),.o(intermediate_reg_1[328]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1472(.clk(clk),.reset(reset),.i1(intermediate_reg_0[655]),.i2(intermediate_reg_0[654]),.o(intermediate_reg_1[327]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1473(.clk(clk),.reset(reset),.i1(intermediate_reg_0[653]),.i2(intermediate_reg_0[652]),.o(intermediate_reg_1[326]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1474(.clk(clk),.reset(reset),.i1(intermediate_reg_0[651]),.i2(intermediate_reg_0[650]),.o(intermediate_reg_1[325])); 
fsm fsm_inst_1_1475(.clk(clk),.reset(reset),.i1(intermediate_reg_0[649]),.i2(intermediate_reg_0[648]),.o(intermediate_reg_1[324])); 
mux_module mux_module_inst_1_1476(.clk(clk),.reset(reset),.i1(intermediate_reg_0[647]),.i2(intermediate_reg_0[646]),.o(intermediate_reg_1[323]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1477(.clk(clk),.reset(reset),.i1(intermediate_reg_0[645]),.i2(intermediate_reg_0[644]),.o(intermediate_reg_1[322])); 
fsm fsm_inst_1_1478(.clk(clk),.reset(reset),.i1(intermediate_reg_0[643]),.i2(intermediate_reg_0[642]),.o(intermediate_reg_1[321])); 
mux_module mux_module_inst_1_1479(.clk(clk),.reset(reset),.i1(intermediate_reg_0[641]),.i2(intermediate_reg_0[640]),.o(intermediate_reg_1[320]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1480(.clk(clk),.reset(reset),.i1(intermediate_reg_0[639]),.i2(intermediate_reg_0[638]),.o(intermediate_reg_1[319])); 
mux_module mux_module_inst_1_1481(.clk(clk),.reset(reset),.i1(intermediate_reg_0[637]),.i2(intermediate_reg_0[636]),.o(intermediate_reg_1[318]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1482(.clk(clk),.reset(reset),.i1(intermediate_reg_0[635]),.i2(intermediate_reg_0[634]),.o(intermediate_reg_1[317]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1483(.clk(clk),.reset(reset),.i1(intermediate_reg_0[633]),.i2(intermediate_reg_0[632]),.o(intermediate_reg_1[316]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1484(.clk(clk),.reset(reset),.i1(intermediate_reg_0[631]),.i2(intermediate_reg_0[630]),.o(intermediate_reg_1[315])); 
mux_module mux_module_inst_1_1485(.clk(clk),.reset(reset),.i1(intermediate_reg_0[629]),.i2(intermediate_reg_0[628]),.o(intermediate_reg_1[314]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1486(.clk(clk),.reset(reset),.i1(intermediate_reg_0[627]),.i2(intermediate_reg_0[626]),.o(intermediate_reg_1[313])); 
fsm fsm_inst_1_1487(.clk(clk),.reset(reset),.i1(intermediate_reg_0[625]),.i2(intermediate_reg_0[624]),.o(intermediate_reg_1[312])); 
fsm fsm_inst_1_1488(.clk(clk),.reset(reset),.i1(intermediate_reg_0[623]),.i2(intermediate_reg_0[622]),.o(intermediate_reg_1[311])); 
mux_module mux_module_inst_1_1489(.clk(clk),.reset(reset),.i1(intermediate_reg_0[621]),.i2(intermediate_reg_0[620]),.o(intermediate_reg_1[310]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1490(.clk(clk),.reset(reset),.i1(intermediate_reg_0[619]),.i2(intermediate_reg_0[618]),.o(intermediate_reg_1[309]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1491(.clk(clk),.reset(reset),.i1(intermediate_reg_0[617]),.i2(intermediate_reg_0[616]),.o(intermediate_reg_1[308]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1492(.clk(clk),.reset(reset),.i1(intermediate_reg_0[615]),.i2(intermediate_reg_0[614]),.o(intermediate_reg_1[307]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1493(.clk(clk),.reset(reset),.i1(intermediate_reg_0[613]),.i2(intermediate_reg_0[612]),.o(intermediate_reg_1[306])); 
mux_module mux_module_inst_1_1494(.clk(clk),.reset(reset),.i1(intermediate_reg_0[611]),.i2(intermediate_reg_0[610]),.o(intermediate_reg_1[305]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1495(.clk(clk),.reset(reset),.i1(intermediate_reg_0[609]),.i2(intermediate_reg_0[608]),.o(intermediate_reg_1[304])); 
fsm fsm_inst_1_1496(.clk(clk),.reset(reset),.i1(intermediate_reg_0[607]),.i2(intermediate_reg_0[606]),.o(intermediate_reg_1[303])); 
fsm fsm_inst_1_1497(.clk(clk),.reset(reset),.i1(intermediate_reg_0[605]),.i2(intermediate_reg_0[604]),.o(intermediate_reg_1[302])); 
fsm fsm_inst_1_1498(.clk(clk),.reset(reset),.i1(intermediate_reg_0[603]),.i2(intermediate_reg_0[602]),.o(intermediate_reg_1[301])); 
fsm fsm_inst_1_1499(.clk(clk),.reset(reset),.i1(intermediate_reg_0[601]),.i2(intermediate_reg_0[600]),.o(intermediate_reg_1[300])); 
mux_module mux_module_inst_1_1500(.clk(clk),.reset(reset),.i1(intermediate_reg_0[599]),.i2(intermediate_reg_0[598]),.o(intermediate_reg_1[299]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1501(.clk(clk),.reset(reset),.i1(intermediate_reg_0[597]),.i2(intermediate_reg_0[596]),.o(intermediate_reg_1[298])); 
mux_module mux_module_inst_1_1502(.clk(clk),.reset(reset),.i1(intermediate_reg_0[595]),.i2(intermediate_reg_0[594]),.o(intermediate_reg_1[297]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1503(.clk(clk),.reset(reset),.i1(intermediate_reg_0[593]),.i2(intermediate_reg_0[592]),.o(intermediate_reg_1[296]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1504(.clk(clk),.reset(reset),.i1(intermediate_reg_0[591]),.i2(intermediate_reg_0[590]),.o(intermediate_reg_1[295]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1505(.clk(clk),.reset(reset),.i1(intermediate_reg_0[589]),.i2(intermediate_reg_0[588]),.o(intermediate_reg_1[294]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1506(.clk(clk),.reset(reset),.i1(intermediate_reg_0[587]),.i2(intermediate_reg_0[586]),.o(intermediate_reg_1[293])); 
fsm fsm_inst_1_1507(.clk(clk),.reset(reset),.i1(intermediate_reg_0[585]),.i2(intermediate_reg_0[584]),.o(intermediate_reg_1[292])); 
mux_module mux_module_inst_1_1508(.clk(clk),.reset(reset),.i1(intermediate_reg_0[583]),.i2(intermediate_reg_0[582]),.o(intermediate_reg_1[291]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1509(.clk(clk),.reset(reset),.i1(intermediate_reg_0[581]),.i2(intermediate_reg_0[580]),.o(intermediate_reg_1[290])); 
mux_module mux_module_inst_1_1510(.clk(clk),.reset(reset),.i1(intermediate_reg_0[579]),.i2(intermediate_reg_0[578]),.o(intermediate_reg_1[289]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1511(.clk(clk),.reset(reset),.i1(intermediate_reg_0[577]),.i2(intermediate_reg_0[576]),.o(intermediate_reg_1[288])); 
fsm fsm_inst_1_1512(.clk(clk),.reset(reset),.i1(intermediate_reg_0[575]),.i2(intermediate_reg_0[574]),.o(intermediate_reg_1[287])); 
fsm fsm_inst_1_1513(.clk(clk),.reset(reset),.i1(intermediate_reg_0[573]),.i2(intermediate_reg_0[572]),.o(intermediate_reg_1[286])); 
fsm fsm_inst_1_1514(.clk(clk),.reset(reset),.i1(intermediate_reg_0[571]),.i2(intermediate_reg_0[570]),.o(intermediate_reg_1[285])); 
mux_module mux_module_inst_1_1515(.clk(clk),.reset(reset),.i1(intermediate_reg_0[569]),.i2(intermediate_reg_0[568]),.o(intermediate_reg_1[284]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1516(.clk(clk),.reset(reset),.i1(intermediate_reg_0[567]),.i2(intermediate_reg_0[566]),.o(intermediate_reg_1[283])); 
fsm fsm_inst_1_1517(.clk(clk),.reset(reset),.i1(intermediate_reg_0[565]),.i2(intermediate_reg_0[564]),.o(intermediate_reg_1[282])); 
fsm fsm_inst_1_1518(.clk(clk),.reset(reset),.i1(intermediate_reg_0[563]),.i2(intermediate_reg_0[562]),.o(intermediate_reg_1[281])); 
mux_module mux_module_inst_1_1519(.clk(clk),.reset(reset),.i1(intermediate_reg_0[561]),.i2(intermediate_reg_0[560]),.o(intermediate_reg_1[280]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1520(.clk(clk),.reset(reset),.i1(intermediate_reg_0[559]),.i2(intermediate_reg_0[558]),.o(intermediate_reg_1[279])); 
mux_module mux_module_inst_1_1521(.clk(clk),.reset(reset),.i1(intermediate_reg_0[557]),.i2(intermediate_reg_0[556]),.o(intermediate_reg_1[278]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1522(.clk(clk),.reset(reset),.i1(intermediate_reg_0[555]),.i2(intermediate_reg_0[554]),.o(intermediate_reg_1[277])); 
fsm fsm_inst_1_1523(.clk(clk),.reset(reset),.i1(intermediate_reg_0[553]),.i2(intermediate_reg_0[552]),.o(intermediate_reg_1[276])); 
fsm fsm_inst_1_1524(.clk(clk),.reset(reset),.i1(intermediate_reg_0[551]),.i2(intermediate_reg_0[550]),.o(intermediate_reg_1[275])); 
fsm fsm_inst_1_1525(.clk(clk),.reset(reset),.i1(intermediate_reg_0[549]),.i2(intermediate_reg_0[548]),.o(intermediate_reg_1[274])); 
fsm fsm_inst_1_1526(.clk(clk),.reset(reset),.i1(intermediate_reg_0[547]),.i2(intermediate_reg_0[546]),.o(intermediate_reg_1[273])); 
fsm fsm_inst_1_1527(.clk(clk),.reset(reset),.i1(intermediate_reg_0[545]),.i2(intermediate_reg_0[544]),.o(intermediate_reg_1[272])); 
mux_module mux_module_inst_1_1528(.clk(clk),.reset(reset),.i1(intermediate_reg_0[543]),.i2(intermediate_reg_0[542]),.o(intermediate_reg_1[271]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1529(.clk(clk),.reset(reset),.i1(intermediate_reg_0[541]),.i2(intermediate_reg_0[540]),.o(intermediate_reg_1[270])); 
fsm fsm_inst_1_1530(.clk(clk),.reset(reset),.i1(intermediate_reg_0[539]),.i2(intermediate_reg_0[538]),.o(intermediate_reg_1[269])); 
fsm fsm_inst_1_1531(.clk(clk),.reset(reset),.i1(intermediate_reg_0[537]),.i2(intermediate_reg_0[536]),.o(intermediate_reg_1[268])); 
fsm fsm_inst_1_1532(.clk(clk),.reset(reset),.i1(intermediate_reg_0[535]),.i2(intermediate_reg_0[534]),.o(intermediate_reg_1[267])); 
fsm fsm_inst_1_1533(.clk(clk),.reset(reset),.i1(intermediate_reg_0[533]),.i2(intermediate_reg_0[532]),.o(intermediate_reg_1[266])); 
fsm fsm_inst_1_1534(.clk(clk),.reset(reset),.i1(intermediate_reg_0[531]),.i2(intermediate_reg_0[530]),.o(intermediate_reg_1[265])); 
mux_module mux_module_inst_1_1535(.clk(clk),.reset(reset),.i1(intermediate_reg_0[529]),.i2(intermediate_reg_0[528]),.o(intermediate_reg_1[264]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1536(.clk(clk),.reset(reset),.i1(intermediate_reg_0[527]),.i2(intermediate_reg_0[526]),.o(intermediate_reg_1[263])); 
fsm fsm_inst_1_1537(.clk(clk),.reset(reset),.i1(intermediate_reg_0[525]),.i2(intermediate_reg_0[524]),.o(intermediate_reg_1[262])); 
fsm fsm_inst_1_1538(.clk(clk),.reset(reset),.i1(intermediate_reg_0[523]),.i2(intermediate_reg_0[522]),.o(intermediate_reg_1[261])); 
fsm fsm_inst_1_1539(.clk(clk),.reset(reset),.i1(intermediate_reg_0[521]),.i2(intermediate_reg_0[520]),.o(intermediate_reg_1[260])); 
mux_module mux_module_inst_1_1540(.clk(clk),.reset(reset),.i1(intermediate_reg_0[519]),.i2(intermediate_reg_0[518]),.o(intermediate_reg_1[259]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1541(.clk(clk),.reset(reset),.i1(intermediate_reg_0[517]),.i2(intermediate_reg_0[516]),.o(intermediate_reg_1[258])); 
mux_module mux_module_inst_1_1542(.clk(clk),.reset(reset),.i1(intermediate_reg_0[515]),.i2(intermediate_reg_0[514]),.o(intermediate_reg_1[257]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1543(.clk(clk),.reset(reset),.i1(intermediate_reg_0[513]),.i2(intermediate_reg_0[512]),.o(intermediate_reg_1[256])); 
mux_module mux_module_inst_1_1544(.clk(clk),.reset(reset),.i1(intermediate_reg_0[511]),.i2(intermediate_reg_0[510]),.o(intermediate_reg_1[255]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1545(.clk(clk),.reset(reset),.i1(intermediate_reg_0[509]),.i2(intermediate_reg_0[508]),.o(intermediate_reg_1[254]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1546(.clk(clk),.reset(reset),.i1(intermediate_reg_0[507]),.i2(intermediate_reg_0[506]),.o(intermediate_reg_1[253])); 
fsm fsm_inst_1_1547(.clk(clk),.reset(reset),.i1(intermediate_reg_0[505]),.i2(intermediate_reg_0[504]),.o(intermediate_reg_1[252])); 
fsm fsm_inst_1_1548(.clk(clk),.reset(reset),.i1(intermediate_reg_0[503]),.i2(intermediate_reg_0[502]),.o(intermediate_reg_1[251])); 
fsm fsm_inst_1_1549(.clk(clk),.reset(reset),.i1(intermediate_reg_0[501]),.i2(intermediate_reg_0[500]),.o(intermediate_reg_1[250])); 
fsm fsm_inst_1_1550(.clk(clk),.reset(reset),.i1(intermediate_reg_0[499]),.i2(intermediate_reg_0[498]),.o(intermediate_reg_1[249])); 
fsm fsm_inst_1_1551(.clk(clk),.reset(reset),.i1(intermediate_reg_0[497]),.i2(intermediate_reg_0[496]),.o(intermediate_reg_1[248])); 
mux_module mux_module_inst_1_1552(.clk(clk),.reset(reset),.i1(intermediate_reg_0[495]),.i2(intermediate_reg_0[494]),.o(intermediate_reg_1[247]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1553(.clk(clk),.reset(reset),.i1(intermediate_reg_0[493]),.i2(intermediate_reg_0[492]),.o(intermediate_reg_1[246]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1554(.clk(clk),.reset(reset),.i1(intermediate_reg_0[491]),.i2(intermediate_reg_0[490]),.o(intermediate_reg_1[245]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1555(.clk(clk),.reset(reset),.i1(intermediate_reg_0[489]),.i2(intermediate_reg_0[488]),.o(intermediate_reg_1[244]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1556(.clk(clk),.reset(reset),.i1(intermediate_reg_0[487]),.i2(intermediate_reg_0[486]),.o(intermediate_reg_1[243])); 
fsm fsm_inst_1_1557(.clk(clk),.reset(reset),.i1(intermediate_reg_0[485]),.i2(intermediate_reg_0[484]),.o(intermediate_reg_1[242])); 
mux_module mux_module_inst_1_1558(.clk(clk),.reset(reset),.i1(intermediate_reg_0[483]),.i2(intermediate_reg_0[482]),.o(intermediate_reg_1[241]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1559(.clk(clk),.reset(reset),.i1(intermediate_reg_0[481]),.i2(intermediate_reg_0[480]),.o(intermediate_reg_1[240])); 
mux_module mux_module_inst_1_1560(.clk(clk),.reset(reset),.i1(intermediate_reg_0[479]),.i2(intermediate_reg_0[478]),.o(intermediate_reg_1[239]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1561(.clk(clk),.reset(reset),.i1(intermediate_reg_0[477]),.i2(intermediate_reg_0[476]),.o(intermediate_reg_1[238]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1562(.clk(clk),.reset(reset),.i1(intermediate_reg_0[475]),.i2(intermediate_reg_0[474]),.o(intermediate_reg_1[237]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1563(.clk(clk),.reset(reset),.i1(intermediate_reg_0[473]),.i2(intermediate_reg_0[472]),.o(intermediate_reg_1[236]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1564(.clk(clk),.reset(reset),.i1(intermediate_reg_0[471]),.i2(intermediate_reg_0[470]),.o(intermediate_reg_1[235]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1565(.clk(clk),.reset(reset),.i1(intermediate_reg_0[469]),.i2(intermediate_reg_0[468]),.o(intermediate_reg_1[234])); 
fsm fsm_inst_1_1566(.clk(clk),.reset(reset),.i1(intermediate_reg_0[467]),.i2(intermediate_reg_0[466]),.o(intermediate_reg_1[233])); 
mux_module mux_module_inst_1_1567(.clk(clk),.reset(reset),.i1(intermediate_reg_0[465]),.i2(intermediate_reg_0[464]),.o(intermediate_reg_1[232]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1568(.clk(clk),.reset(reset),.i1(intermediate_reg_0[463]),.i2(intermediate_reg_0[462]),.o(intermediate_reg_1[231])); 
fsm fsm_inst_1_1569(.clk(clk),.reset(reset),.i1(intermediate_reg_0[461]),.i2(intermediate_reg_0[460]),.o(intermediate_reg_1[230])); 
mux_module mux_module_inst_1_1570(.clk(clk),.reset(reset),.i1(intermediate_reg_0[459]),.i2(intermediate_reg_0[458]),.o(intermediate_reg_1[229]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1571(.clk(clk),.reset(reset),.i1(intermediate_reg_0[457]),.i2(intermediate_reg_0[456]),.o(intermediate_reg_1[228])); 
fsm fsm_inst_1_1572(.clk(clk),.reset(reset),.i1(intermediate_reg_0[455]),.i2(intermediate_reg_0[454]),.o(intermediate_reg_1[227])); 
fsm fsm_inst_1_1573(.clk(clk),.reset(reset),.i1(intermediate_reg_0[453]),.i2(intermediate_reg_0[452]),.o(intermediate_reg_1[226])); 
mux_module mux_module_inst_1_1574(.clk(clk),.reset(reset),.i1(intermediate_reg_0[451]),.i2(intermediate_reg_0[450]),.o(intermediate_reg_1[225]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1575(.clk(clk),.reset(reset),.i1(intermediate_reg_0[449]),.i2(intermediate_reg_0[448]),.o(intermediate_reg_1[224])); 
fsm fsm_inst_1_1576(.clk(clk),.reset(reset),.i1(intermediate_reg_0[447]),.i2(intermediate_reg_0[446]),.o(intermediate_reg_1[223])); 
mux_module mux_module_inst_1_1577(.clk(clk),.reset(reset),.i1(intermediate_reg_0[445]),.i2(intermediate_reg_0[444]),.o(intermediate_reg_1[222]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1578(.clk(clk),.reset(reset),.i1(intermediate_reg_0[443]),.i2(intermediate_reg_0[442]),.o(intermediate_reg_1[221]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1579(.clk(clk),.reset(reset),.i1(intermediate_reg_0[441]),.i2(intermediate_reg_0[440]),.o(intermediate_reg_1[220])); 
mux_module mux_module_inst_1_1580(.clk(clk),.reset(reset),.i1(intermediate_reg_0[439]),.i2(intermediate_reg_0[438]),.o(intermediate_reg_1[219]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1581(.clk(clk),.reset(reset),.i1(intermediate_reg_0[437]),.i2(intermediate_reg_0[436]),.o(intermediate_reg_1[218]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1582(.clk(clk),.reset(reset),.i1(intermediate_reg_0[435]),.i2(intermediate_reg_0[434]),.o(intermediate_reg_1[217]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1583(.clk(clk),.reset(reset),.i1(intermediate_reg_0[433]),.i2(intermediate_reg_0[432]),.o(intermediate_reg_1[216]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1584(.clk(clk),.reset(reset),.i1(intermediate_reg_0[431]),.i2(intermediate_reg_0[430]),.o(intermediate_reg_1[215])); 
mux_module mux_module_inst_1_1585(.clk(clk),.reset(reset),.i1(intermediate_reg_0[429]),.i2(intermediate_reg_0[428]),.o(intermediate_reg_1[214]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1586(.clk(clk),.reset(reset),.i1(intermediate_reg_0[427]),.i2(intermediate_reg_0[426]),.o(intermediate_reg_1[213]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1587(.clk(clk),.reset(reset),.i1(intermediate_reg_0[425]),.i2(intermediate_reg_0[424]),.o(intermediate_reg_1[212])); 
fsm fsm_inst_1_1588(.clk(clk),.reset(reset),.i1(intermediate_reg_0[423]),.i2(intermediate_reg_0[422]),.o(intermediate_reg_1[211])); 
fsm fsm_inst_1_1589(.clk(clk),.reset(reset),.i1(intermediate_reg_0[421]),.i2(intermediate_reg_0[420]),.o(intermediate_reg_1[210])); 
mux_module mux_module_inst_1_1590(.clk(clk),.reset(reset),.i1(intermediate_reg_0[419]),.i2(intermediate_reg_0[418]),.o(intermediate_reg_1[209]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1591(.clk(clk),.reset(reset),.i1(intermediate_reg_0[417]),.i2(intermediate_reg_0[416]),.o(intermediate_reg_1[208])); 
fsm fsm_inst_1_1592(.clk(clk),.reset(reset),.i1(intermediate_reg_0[415]),.i2(intermediate_reg_0[414]),.o(intermediate_reg_1[207])); 
mux_module mux_module_inst_1_1593(.clk(clk),.reset(reset),.i1(intermediate_reg_0[413]),.i2(intermediate_reg_0[412]),.o(intermediate_reg_1[206]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1594(.clk(clk),.reset(reset),.i1(intermediate_reg_0[411]),.i2(intermediate_reg_0[410]),.o(intermediate_reg_1[205])); 
fsm fsm_inst_1_1595(.clk(clk),.reset(reset),.i1(intermediate_reg_0[409]),.i2(intermediate_reg_0[408]),.o(intermediate_reg_1[204])); 
fsm fsm_inst_1_1596(.clk(clk),.reset(reset),.i1(intermediate_reg_0[407]),.i2(intermediate_reg_0[406]),.o(intermediate_reg_1[203])); 
fsm fsm_inst_1_1597(.clk(clk),.reset(reset),.i1(intermediate_reg_0[405]),.i2(intermediate_reg_0[404]),.o(intermediate_reg_1[202])); 
fsm fsm_inst_1_1598(.clk(clk),.reset(reset),.i1(intermediate_reg_0[403]),.i2(intermediate_reg_0[402]),.o(intermediate_reg_1[201])); 
mux_module mux_module_inst_1_1599(.clk(clk),.reset(reset),.i1(intermediate_reg_0[401]),.i2(intermediate_reg_0[400]),.o(intermediate_reg_1[200]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1600(.clk(clk),.reset(reset),.i1(intermediate_reg_0[399]),.i2(intermediate_reg_0[398]),.o(intermediate_reg_1[199]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1601(.clk(clk),.reset(reset),.i1(intermediate_reg_0[397]),.i2(intermediate_reg_0[396]),.o(intermediate_reg_1[198])); 
fsm fsm_inst_1_1602(.clk(clk),.reset(reset),.i1(intermediate_reg_0[395]),.i2(intermediate_reg_0[394]),.o(intermediate_reg_1[197])); 
mux_module mux_module_inst_1_1603(.clk(clk),.reset(reset),.i1(intermediate_reg_0[393]),.i2(intermediate_reg_0[392]),.o(intermediate_reg_1[196]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1604(.clk(clk),.reset(reset),.i1(intermediate_reg_0[391]),.i2(intermediate_reg_0[390]),.o(intermediate_reg_1[195]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1605(.clk(clk),.reset(reset),.i1(intermediate_reg_0[389]),.i2(intermediate_reg_0[388]),.o(intermediate_reg_1[194]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1606(.clk(clk),.reset(reset),.i1(intermediate_reg_0[387]),.i2(intermediate_reg_0[386]),.o(intermediate_reg_1[193]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1607(.clk(clk),.reset(reset),.i1(intermediate_reg_0[385]),.i2(intermediate_reg_0[384]),.o(intermediate_reg_1[192])); 
mux_module mux_module_inst_1_1608(.clk(clk),.reset(reset),.i1(intermediate_reg_0[383]),.i2(intermediate_reg_0[382]),.o(intermediate_reg_1[191]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1609(.clk(clk),.reset(reset),.i1(intermediate_reg_0[381]),.i2(intermediate_reg_0[380]),.o(intermediate_reg_1[190])); 
fsm fsm_inst_1_1610(.clk(clk),.reset(reset),.i1(intermediate_reg_0[379]),.i2(intermediate_reg_0[378]),.o(intermediate_reg_1[189])); 
fsm fsm_inst_1_1611(.clk(clk),.reset(reset),.i1(intermediate_reg_0[377]),.i2(intermediate_reg_0[376]),.o(intermediate_reg_1[188])); 
fsm fsm_inst_1_1612(.clk(clk),.reset(reset),.i1(intermediate_reg_0[375]),.i2(intermediate_reg_0[374]),.o(intermediate_reg_1[187])); 
fsm fsm_inst_1_1613(.clk(clk),.reset(reset),.i1(intermediate_reg_0[373]),.i2(intermediate_reg_0[372]),.o(intermediate_reg_1[186])); 
mux_module mux_module_inst_1_1614(.clk(clk),.reset(reset),.i1(intermediate_reg_0[371]),.i2(intermediate_reg_0[370]),.o(intermediate_reg_1[185]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1615(.clk(clk),.reset(reset),.i1(intermediate_reg_0[369]),.i2(intermediate_reg_0[368]),.o(intermediate_reg_1[184])); 
fsm fsm_inst_1_1616(.clk(clk),.reset(reset),.i1(intermediate_reg_0[367]),.i2(intermediate_reg_0[366]),.o(intermediate_reg_1[183])); 
fsm fsm_inst_1_1617(.clk(clk),.reset(reset),.i1(intermediate_reg_0[365]),.i2(intermediate_reg_0[364]),.o(intermediate_reg_1[182])); 
mux_module mux_module_inst_1_1618(.clk(clk),.reset(reset),.i1(intermediate_reg_0[363]),.i2(intermediate_reg_0[362]),.o(intermediate_reg_1[181]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1619(.clk(clk),.reset(reset),.i1(intermediate_reg_0[361]),.i2(intermediate_reg_0[360]),.o(intermediate_reg_1[180]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1620(.clk(clk),.reset(reset),.i1(intermediate_reg_0[359]),.i2(intermediate_reg_0[358]),.o(intermediate_reg_1[179])); 
fsm fsm_inst_1_1621(.clk(clk),.reset(reset),.i1(intermediate_reg_0[357]),.i2(intermediate_reg_0[356]),.o(intermediate_reg_1[178])); 
mux_module mux_module_inst_1_1622(.clk(clk),.reset(reset),.i1(intermediate_reg_0[355]),.i2(intermediate_reg_0[354]),.o(intermediate_reg_1[177]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1623(.clk(clk),.reset(reset),.i1(intermediate_reg_0[353]),.i2(intermediate_reg_0[352]),.o(intermediate_reg_1[176])); 
fsm fsm_inst_1_1624(.clk(clk),.reset(reset),.i1(intermediate_reg_0[351]),.i2(intermediate_reg_0[350]),.o(intermediate_reg_1[175])); 
mux_module mux_module_inst_1_1625(.clk(clk),.reset(reset),.i1(intermediate_reg_0[349]),.i2(intermediate_reg_0[348]),.o(intermediate_reg_1[174]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1626(.clk(clk),.reset(reset),.i1(intermediate_reg_0[347]),.i2(intermediate_reg_0[346]),.o(intermediate_reg_1[173])); 
fsm fsm_inst_1_1627(.clk(clk),.reset(reset),.i1(intermediate_reg_0[345]),.i2(intermediate_reg_0[344]),.o(intermediate_reg_1[172])); 
fsm fsm_inst_1_1628(.clk(clk),.reset(reset),.i1(intermediate_reg_0[343]),.i2(intermediate_reg_0[342]),.o(intermediate_reg_1[171])); 
mux_module mux_module_inst_1_1629(.clk(clk),.reset(reset),.i1(intermediate_reg_0[341]),.i2(intermediate_reg_0[340]),.o(intermediate_reg_1[170]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1630(.clk(clk),.reset(reset),.i1(intermediate_reg_0[339]),.i2(intermediate_reg_0[338]),.o(intermediate_reg_1[169]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1631(.clk(clk),.reset(reset),.i1(intermediate_reg_0[337]),.i2(intermediate_reg_0[336]),.o(intermediate_reg_1[168]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1632(.clk(clk),.reset(reset),.i1(intermediate_reg_0[335]),.i2(intermediate_reg_0[334]),.o(intermediate_reg_1[167]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1633(.clk(clk),.reset(reset),.i1(intermediate_reg_0[333]),.i2(intermediate_reg_0[332]),.o(intermediate_reg_1[166]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1634(.clk(clk),.reset(reset),.i1(intermediate_reg_0[331]),.i2(intermediate_reg_0[330]),.o(intermediate_reg_1[165])); 
fsm fsm_inst_1_1635(.clk(clk),.reset(reset),.i1(intermediate_reg_0[329]),.i2(intermediate_reg_0[328]),.o(intermediate_reg_1[164])); 
fsm fsm_inst_1_1636(.clk(clk),.reset(reset),.i1(intermediate_reg_0[327]),.i2(intermediate_reg_0[326]),.o(intermediate_reg_1[163])); 
fsm fsm_inst_1_1637(.clk(clk),.reset(reset),.i1(intermediate_reg_0[325]),.i2(intermediate_reg_0[324]),.o(intermediate_reg_1[162])); 
mux_module mux_module_inst_1_1638(.clk(clk),.reset(reset),.i1(intermediate_reg_0[323]),.i2(intermediate_reg_0[322]),.o(intermediate_reg_1[161]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1639(.clk(clk),.reset(reset),.i1(intermediate_reg_0[321]),.i2(intermediate_reg_0[320]),.o(intermediate_reg_1[160])); 
mux_module mux_module_inst_1_1640(.clk(clk),.reset(reset),.i1(intermediate_reg_0[319]),.i2(intermediate_reg_0[318]),.o(intermediate_reg_1[159]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1641(.clk(clk),.reset(reset),.i1(intermediate_reg_0[317]),.i2(intermediate_reg_0[316]),.o(intermediate_reg_1[158]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1642(.clk(clk),.reset(reset),.i1(intermediate_reg_0[315]),.i2(intermediate_reg_0[314]),.o(intermediate_reg_1[157]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1643(.clk(clk),.reset(reset),.i1(intermediate_reg_0[313]),.i2(intermediate_reg_0[312]),.o(intermediate_reg_1[156])); 
mux_module mux_module_inst_1_1644(.clk(clk),.reset(reset),.i1(intermediate_reg_0[311]),.i2(intermediate_reg_0[310]),.o(intermediate_reg_1[155]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1645(.clk(clk),.reset(reset),.i1(intermediate_reg_0[309]),.i2(intermediate_reg_0[308]),.o(intermediate_reg_1[154])); 
fsm fsm_inst_1_1646(.clk(clk),.reset(reset),.i1(intermediate_reg_0[307]),.i2(intermediate_reg_0[306]),.o(intermediate_reg_1[153])); 
mux_module mux_module_inst_1_1647(.clk(clk),.reset(reset),.i1(intermediate_reg_0[305]),.i2(intermediate_reg_0[304]),.o(intermediate_reg_1[152]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1648(.clk(clk),.reset(reset),.i1(intermediate_reg_0[303]),.i2(intermediate_reg_0[302]),.o(intermediate_reg_1[151])); 
mux_module mux_module_inst_1_1649(.clk(clk),.reset(reset),.i1(intermediate_reg_0[301]),.i2(intermediate_reg_0[300]),.o(intermediate_reg_1[150]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1650(.clk(clk),.reset(reset),.i1(intermediate_reg_0[299]),.i2(intermediate_reg_0[298]),.o(intermediate_reg_1[149])); 
mux_module mux_module_inst_1_1651(.clk(clk),.reset(reset),.i1(intermediate_reg_0[297]),.i2(intermediate_reg_0[296]),.o(intermediate_reg_1[148]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1652(.clk(clk),.reset(reset),.i1(intermediate_reg_0[295]),.i2(intermediate_reg_0[294]),.o(intermediate_reg_1[147])); 
mux_module mux_module_inst_1_1653(.clk(clk),.reset(reset),.i1(intermediate_reg_0[293]),.i2(intermediate_reg_0[292]),.o(intermediate_reg_1[146]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1654(.clk(clk),.reset(reset),.i1(intermediate_reg_0[291]),.i2(intermediate_reg_0[290]),.o(intermediate_reg_1[145])); 
fsm fsm_inst_1_1655(.clk(clk),.reset(reset),.i1(intermediate_reg_0[289]),.i2(intermediate_reg_0[288]),.o(intermediate_reg_1[144])); 
fsm fsm_inst_1_1656(.clk(clk),.reset(reset),.i1(intermediate_reg_0[287]),.i2(intermediate_reg_0[286]),.o(intermediate_reg_1[143])); 
fsm fsm_inst_1_1657(.clk(clk),.reset(reset),.i1(intermediate_reg_0[285]),.i2(intermediate_reg_0[284]),.o(intermediate_reg_1[142])); 
fsm fsm_inst_1_1658(.clk(clk),.reset(reset),.i1(intermediate_reg_0[283]),.i2(intermediate_reg_0[282]),.o(intermediate_reg_1[141])); 
fsm fsm_inst_1_1659(.clk(clk),.reset(reset),.i1(intermediate_reg_0[281]),.i2(intermediate_reg_0[280]),.o(intermediate_reg_1[140])); 
mux_module mux_module_inst_1_1660(.clk(clk),.reset(reset),.i1(intermediate_reg_0[279]),.i2(intermediate_reg_0[278]),.o(intermediate_reg_1[139]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1661(.clk(clk),.reset(reset),.i1(intermediate_reg_0[277]),.i2(intermediate_reg_0[276]),.o(intermediate_reg_1[138]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1662(.clk(clk),.reset(reset),.i1(intermediate_reg_0[275]),.i2(intermediate_reg_0[274]),.o(intermediate_reg_1[137]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1663(.clk(clk),.reset(reset),.i1(intermediate_reg_0[273]),.i2(intermediate_reg_0[272]),.o(intermediate_reg_1[136])); 
fsm fsm_inst_1_1664(.clk(clk),.reset(reset),.i1(intermediate_reg_0[271]),.i2(intermediate_reg_0[270]),.o(intermediate_reg_1[135])); 
fsm fsm_inst_1_1665(.clk(clk),.reset(reset),.i1(intermediate_reg_0[269]),.i2(intermediate_reg_0[268]),.o(intermediate_reg_1[134])); 
fsm fsm_inst_1_1666(.clk(clk),.reset(reset),.i1(intermediate_reg_0[267]),.i2(intermediate_reg_0[266]),.o(intermediate_reg_1[133])); 
fsm fsm_inst_1_1667(.clk(clk),.reset(reset),.i1(intermediate_reg_0[265]),.i2(intermediate_reg_0[264]),.o(intermediate_reg_1[132])); 
fsm fsm_inst_1_1668(.clk(clk),.reset(reset),.i1(intermediate_reg_0[263]),.i2(intermediate_reg_0[262]),.o(intermediate_reg_1[131])); 
fsm fsm_inst_1_1669(.clk(clk),.reset(reset),.i1(intermediate_reg_0[261]),.i2(intermediate_reg_0[260]),.o(intermediate_reg_1[130])); 
mux_module mux_module_inst_1_1670(.clk(clk),.reset(reset),.i1(intermediate_reg_0[259]),.i2(intermediate_reg_0[258]),.o(intermediate_reg_1[129]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1671(.clk(clk),.reset(reset),.i1(intermediate_reg_0[257]),.i2(intermediate_reg_0[256]),.o(intermediate_reg_1[128])); 
mux_module mux_module_inst_1_1672(.clk(clk),.reset(reset),.i1(intermediate_reg_0[255]),.i2(intermediate_reg_0[254]),.o(intermediate_reg_1[127]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1673(.clk(clk),.reset(reset),.i1(intermediate_reg_0[253]),.i2(intermediate_reg_0[252]),.o(intermediate_reg_1[126])); 
mux_module mux_module_inst_1_1674(.clk(clk),.reset(reset),.i1(intermediate_reg_0[251]),.i2(intermediate_reg_0[250]),.o(intermediate_reg_1[125]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1675(.clk(clk),.reset(reset),.i1(intermediate_reg_0[249]),.i2(intermediate_reg_0[248]),.o(intermediate_reg_1[124])); 
mux_module mux_module_inst_1_1676(.clk(clk),.reset(reset),.i1(intermediate_reg_0[247]),.i2(intermediate_reg_0[246]),.o(intermediate_reg_1[123]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1677(.clk(clk),.reset(reset),.i1(intermediate_reg_0[245]),.i2(intermediate_reg_0[244]),.o(intermediate_reg_1[122])); 
mux_module mux_module_inst_1_1678(.clk(clk),.reset(reset),.i1(intermediate_reg_0[243]),.i2(intermediate_reg_0[242]),.o(intermediate_reg_1[121]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1679(.clk(clk),.reset(reset),.i1(intermediate_reg_0[241]),.i2(intermediate_reg_0[240]),.o(intermediate_reg_1[120])); 
mux_module mux_module_inst_1_1680(.clk(clk),.reset(reset),.i1(intermediate_reg_0[239]),.i2(intermediate_reg_0[238]),.o(intermediate_reg_1[119]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1681(.clk(clk),.reset(reset),.i1(intermediate_reg_0[237]),.i2(intermediate_reg_0[236]),.o(intermediate_reg_1[118]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1682(.clk(clk),.reset(reset),.i1(intermediate_reg_0[235]),.i2(intermediate_reg_0[234]),.o(intermediate_reg_1[117]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1683(.clk(clk),.reset(reset),.i1(intermediate_reg_0[233]),.i2(intermediate_reg_0[232]),.o(intermediate_reg_1[116]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1684(.clk(clk),.reset(reset),.i1(intermediate_reg_0[231]),.i2(intermediate_reg_0[230]),.o(intermediate_reg_1[115]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1685(.clk(clk),.reset(reset),.i1(intermediate_reg_0[229]),.i2(intermediate_reg_0[228]),.o(intermediate_reg_1[114])); 
mux_module mux_module_inst_1_1686(.clk(clk),.reset(reset),.i1(intermediate_reg_0[227]),.i2(intermediate_reg_0[226]),.o(intermediate_reg_1[113]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1687(.clk(clk),.reset(reset),.i1(intermediate_reg_0[225]),.i2(intermediate_reg_0[224]),.o(intermediate_reg_1[112]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1688(.clk(clk),.reset(reset),.i1(intermediate_reg_0[223]),.i2(intermediate_reg_0[222]),.o(intermediate_reg_1[111]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1689(.clk(clk),.reset(reset),.i1(intermediate_reg_0[221]),.i2(intermediate_reg_0[220]),.o(intermediate_reg_1[110])); 
mux_module mux_module_inst_1_1690(.clk(clk),.reset(reset),.i1(intermediate_reg_0[219]),.i2(intermediate_reg_0[218]),.o(intermediate_reg_1[109]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1691(.clk(clk),.reset(reset),.i1(intermediate_reg_0[217]),.i2(intermediate_reg_0[216]),.o(intermediate_reg_1[108]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1692(.clk(clk),.reset(reset),.i1(intermediate_reg_0[215]),.i2(intermediate_reg_0[214]),.o(intermediate_reg_1[107]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1693(.clk(clk),.reset(reset),.i1(intermediate_reg_0[213]),.i2(intermediate_reg_0[212]),.o(intermediate_reg_1[106]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1694(.clk(clk),.reset(reset),.i1(intermediate_reg_0[211]),.i2(intermediate_reg_0[210]),.o(intermediate_reg_1[105])); 
mux_module mux_module_inst_1_1695(.clk(clk),.reset(reset),.i1(intermediate_reg_0[209]),.i2(intermediate_reg_0[208]),.o(intermediate_reg_1[104]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1696(.clk(clk),.reset(reset),.i1(intermediate_reg_0[207]),.i2(intermediate_reg_0[206]),.o(intermediate_reg_1[103])); 
mux_module mux_module_inst_1_1697(.clk(clk),.reset(reset),.i1(intermediate_reg_0[205]),.i2(intermediate_reg_0[204]),.o(intermediate_reg_1[102]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1698(.clk(clk),.reset(reset),.i1(intermediate_reg_0[203]),.i2(intermediate_reg_0[202]),.o(intermediate_reg_1[101]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1699(.clk(clk),.reset(reset),.i1(intermediate_reg_0[201]),.i2(intermediate_reg_0[200]),.o(intermediate_reg_1[100]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1700(.clk(clk),.reset(reset),.i1(intermediate_reg_0[199]),.i2(intermediate_reg_0[198]),.o(intermediate_reg_1[99]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1701(.clk(clk),.reset(reset),.i1(intermediate_reg_0[197]),.i2(intermediate_reg_0[196]),.o(intermediate_reg_1[98])); 
fsm fsm_inst_1_1702(.clk(clk),.reset(reset),.i1(intermediate_reg_0[195]),.i2(intermediate_reg_0[194]),.o(intermediate_reg_1[97])); 
mux_module mux_module_inst_1_1703(.clk(clk),.reset(reset),.i1(intermediate_reg_0[193]),.i2(intermediate_reg_0[192]),.o(intermediate_reg_1[96]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1704(.clk(clk),.reset(reset),.i1(intermediate_reg_0[191]),.i2(intermediate_reg_0[190]),.o(intermediate_reg_1[95]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1705(.clk(clk),.reset(reset),.i1(intermediate_reg_0[189]),.i2(intermediate_reg_0[188]),.o(intermediate_reg_1[94]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1706(.clk(clk),.reset(reset),.i1(intermediate_reg_0[187]),.i2(intermediate_reg_0[186]),.o(intermediate_reg_1[93]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1707(.clk(clk),.reset(reset),.i1(intermediate_reg_0[185]),.i2(intermediate_reg_0[184]),.o(intermediate_reg_1[92])); 
mux_module mux_module_inst_1_1708(.clk(clk),.reset(reset),.i1(intermediate_reg_0[183]),.i2(intermediate_reg_0[182]),.o(intermediate_reg_1[91]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1709(.clk(clk),.reset(reset),.i1(intermediate_reg_0[181]),.i2(intermediate_reg_0[180]),.o(intermediate_reg_1[90]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1710(.clk(clk),.reset(reset),.i1(intermediate_reg_0[179]),.i2(intermediate_reg_0[178]),.o(intermediate_reg_1[89]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1711(.clk(clk),.reset(reset),.i1(intermediate_reg_0[177]),.i2(intermediate_reg_0[176]),.o(intermediate_reg_1[88]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1712(.clk(clk),.reset(reset),.i1(intermediate_reg_0[175]),.i2(intermediate_reg_0[174]),.o(intermediate_reg_1[87]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1713(.clk(clk),.reset(reset),.i1(intermediate_reg_0[173]),.i2(intermediate_reg_0[172]),.o(intermediate_reg_1[86]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1714(.clk(clk),.reset(reset),.i1(intermediate_reg_0[171]),.i2(intermediate_reg_0[170]),.o(intermediate_reg_1[85])); 
fsm fsm_inst_1_1715(.clk(clk),.reset(reset),.i1(intermediate_reg_0[169]),.i2(intermediate_reg_0[168]),.o(intermediate_reg_1[84])); 
fsm fsm_inst_1_1716(.clk(clk),.reset(reset),.i1(intermediate_reg_0[167]),.i2(intermediate_reg_0[166]),.o(intermediate_reg_1[83])); 
mux_module mux_module_inst_1_1717(.clk(clk),.reset(reset),.i1(intermediate_reg_0[165]),.i2(intermediate_reg_0[164]),.o(intermediate_reg_1[82]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1718(.clk(clk),.reset(reset),.i1(intermediate_reg_0[163]),.i2(intermediate_reg_0[162]),.o(intermediate_reg_1[81])); 
mux_module mux_module_inst_1_1719(.clk(clk),.reset(reset),.i1(intermediate_reg_0[161]),.i2(intermediate_reg_0[160]),.o(intermediate_reg_1[80]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1720(.clk(clk),.reset(reset),.i1(intermediate_reg_0[159]),.i2(intermediate_reg_0[158]),.o(intermediate_reg_1[79])); 
mux_module mux_module_inst_1_1721(.clk(clk),.reset(reset),.i1(intermediate_reg_0[157]),.i2(intermediate_reg_0[156]),.o(intermediate_reg_1[78]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1722(.clk(clk),.reset(reset),.i1(intermediate_reg_0[155]),.i2(intermediate_reg_0[154]),.o(intermediate_reg_1[77]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1723(.clk(clk),.reset(reset),.i1(intermediate_reg_0[153]),.i2(intermediate_reg_0[152]),.o(intermediate_reg_1[76]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1724(.clk(clk),.reset(reset),.i1(intermediate_reg_0[151]),.i2(intermediate_reg_0[150]),.o(intermediate_reg_1[75]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1725(.clk(clk),.reset(reset),.i1(intermediate_reg_0[149]),.i2(intermediate_reg_0[148]),.o(intermediate_reg_1[74]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1726(.clk(clk),.reset(reset),.i1(intermediate_reg_0[147]),.i2(intermediate_reg_0[146]),.o(intermediate_reg_1[73]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1727(.clk(clk),.reset(reset),.i1(intermediate_reg_0[145]),.i2(intermediate_reg_0[144]),.o(intermediate_reg_1[72])); 
mux_module mux_module_inst_1_1728(.clk(clk),.reset(reset),.i1(intermediate_reg_0[143]),.i2(intermediate_reg_0[142]),.o(intermediate_reg_1[71]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1729(.clk(clk),.reset(reset),.i1(intermediate_reg_0[141]),.i2(intermediate_reg_0[140]),.o(intermediate_reg_1[70])); 
fsm fsm_inst_1_1730(.clk(clk),.reset(reset),.i1(intermediate_reg_0[139]),.i2(intermediate_reg_0[138]),.o(intermediate_reg_1[69])); 
mux_module mux_module_inst_1_1731(.clk(clk),.reset(reset),.i1(intermediate_reg_0[137]),.i2(intermediate_reg_0[136]),.o(intermediate_reg_1[68]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1732(.clk(clk),.reset(reset),.i1(intermediate_reg_0[135]),.i2(intermediate_reg_0[134]),.o(intermediate_reg_1[67])); 
fsm fsm_inst_1_1733(.clk(clk),.reset(reset),.i1(intermediate_reg_0[133]),.i2(intermediate_reg_0[132]),.o(intermediate_reg_1[66])); 
mux_module mux_module_inst_1_1734(.clk(clk),.reset(reset),.i1(intermediate_reg_0[131]),.i2(intermediate_reg_0[130]),.o(intermediate_reg_1[65]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1735(.clk(clk),.reset(reset),.i1(intermediate_reg_0[129]),.i2(intermediate_reg_0[128]),.o(intermediate_reg_1[64]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1736(.clk(clk),.reset(reset),.i1(intermediate_reg_0[127]),.i2(intermediate_reg_0[126]),.o(intermediate_reg_1[63])); 
mux_module mux_module_inst_1_1737(.clk(clk),.reset(reset),.i1(intermediate_reg_0[125]),.i2(intermediate_reg_0[124]),.o(intermediate_reg_1[62]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1738(.clk(clk),.reset(reset),.i1(intermediate_reg_0[123]),.i2(intermediate_reg_0[122]),.o(intermediate_reg_1[61])); 
mux_module mux_module_inst_1_1739(.clk(clk),.reset(reset),.i1(intermediate_reg_0[121]),.i2(intermediate_reg_0[120]),.o(intermediate_reg_1[60]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1740(.clk(clk),.reset(reset),.i1(intermediate_reg_0[119]),.i2(intermediate_reg_0[118]),.o(intermediate_reg_1[59])); 
mux_module mux_module_inst_1_1741(.clk(clk),.reset(reset),.i1(intermediate_reg_0[117]),.i2(intermediate_reg_0[116]),.o(intermediate_reg_1[58]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1742(.clk(clk),.reset(reset),.i1(intermediate_reg_0[115]),.i2(intermediate_reg_0[114]),.o(intermediate_reg_1[57]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1743(.clk(clk),.reset(reset),.i1(intermediate_reg_0[113]),.i2(intermediate_reg_0[112]),.o(intermediate_reg_1[56]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1744(.clk(clk),.reset(reset),.i1(intermediate_reg_0[111]),.i2(intermediate_reg_0[110]),.o(intermediate_reg_1[55])); 
mux_module mux_module_inst_1_1745(.clk(clk),.reset(reset),.i1(intermediate_reg_0[109]),.i2(intermediate_reg_0[108]),.o(intermediate_reg_1[54]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1746(.clk(clk),.reset(reset),.i1(intermediate_reg_0[107]),.i2(intermediate_reg_0[106]),.o(intermediate_reg_1[53]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1747(.clk(clk),.reset(reset),.i1(intermediate_reg_0[105]),.i2(intermediate_reg_0[104]),.o(intermediate_reg_1[52]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1748(.clk(clk),.reset(reset),.i1(intermediate_reg_0[103]),.i2(intermediate_reg_0[102]),.o(intermediate_reg_1[51]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1749(.clk(clk),.reset(reset),.i1(intermediate_reg_0[101]),.i2(intermediate_reg_0[100]),.o(intermediate_reg_1[50])); 
fsm fsm_inst_1_1750(.clk(clk),.reset(reset),.i1(intermediate_reg_0[99]),.i2(intermediate_reg_0[98]),.o(intermediate_reg_1[49])); 
mux_module mux_module_inst_1_1751(.clk(clk),.reset(reset),.i1(intermediate_reg_0[97]),.i2(intermediate_reg_0[96]),.o(intermediate_reg_1[48]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1752(.clk(clk),.reset(reset),.i1(intermediate_reg_0[95]),.i2(intermediate_reg_0[94]),.o(intermediate_reg_1[47])); 
fsm fsm_inst_1_1753(.clk(clk),.reset(reset),.i1(intermediate_reg_0[93]),.i2(intermediate_reg_0[92]),.o(intermediate_reg_1[46])); 
fsm fsm_inst_1_1754(.clk(clk),.reset(reset),.i1(intermediate_reg_0[91]),.i2(intermediate_reg_0[90]),.o(intermediate_reg_1[45])); 
fsm fsm_inst_1_1755(.clk(clk),.reset(reset),.i1(intermediate_reg_0[89]),.i2(intermediate_reg_0[88]),.o(intermediate_reg_1[44])); 
mux_module mux_module_inst_1_1756(.clk(clk),.reset(reset),.i1(intermediate_reg_0[87]),.i2(intermediate_reg_0[86]),.o(intermediate_reg_1[43]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1757(.clk(clk),.reset(reset),.i1(intermediate_reg_0[85]),.i2(intermediate_reg_0[84]),.o(intermediate_reg_1[42])); 
fsm fsm_inst_1_1758(.clk(clk),.reset(reset),.i1(intermediate_reg_0[83]),.i2(intermediate_reg_0[82]),.o(intermediate_reg_1[41])); 
fsm fsm_inst_1_1759(.clk(clk),.reset(reset),.i1(intermediate_reg_0[81]),.i2(intermediate_reg_0[80]),.o(intermediate_reg_1[40])); 
mux_module mux_module_inst_1_1760(.clk(clk),.reset(reset),.i1(intermediate_reg_0[79]),.i2(intermediate_reg_0[78]),.o(intermediate_reg_1[39]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1761(.clk(clk),.reset(reset),.i1(intermediate_reg_0[77]),.i2(intermediate_reg_0[76]),.o(intermediate_reg_1[38]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1762(.clk(clk),.reset(reset),.i1(intermediate_reg_0[75]),.i2(intermediate_reg_0[74]),.o(intermediate_reg_1[37]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1763(.clk(clk),.reset(reset),.i1(intermediate_reg_0[73]),.i2(intermediate_reg_0[72]),.o(intermediate_reg_1[36]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1764(.clk(clk),.reset(reset),.i1(intermediate_reg_0[71]),.i2(intermediate_reg_0[70]),.o(intermediate_reg_1[35]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1765(.clk(clk),.reset(reset),.i1(intermediate_reg_0[69]),.i2(intermediate_reg_0[68]),.o(intermediate_reg_1[34])); 
fsm fsm_inst_1_1766(.clk(clk),.reset(reset),.i1(intermediate_reg_0[67]),.i2(intermediate_reg_0[66]),.o(intermediate_reg_1[33])); 
mux_module mux_module_inst_1_1767(.clk(clk),.reset(reset),.i1(intermediate_reg_0[65]),.i2(intermediate_reg_0[64]),.o(intermediate_reg_1[32]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1768(.clk(clk),.reset(reset),.i1(intermediate_reg_0[63]),.i2(intermediate_reg_0[62]),.o(intermediate_reg_1[31])); 
mux_module mux_module_inst_1_1769(.clk(clk),.reset(reset),.i1(intermediate_reg_0[61]),.i2(intermediate_reg_0[60]),.o(intermediate_reg_1[30]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1770(.clk(clk),.reset(reset),.i1(intermediate_reg_0[59]),.i2(intermediate_reg_0[58]),.o(intermediate_reg_1[29])); 
fsm fsm_inst_1_1771(.clk(clk),.reset(reset),.i1(intermediate_reg_0[57]),.i2(intermediate_reg_0[56]),.o(intermediate_reg_1[28])); 
mux_module mux_module_inst_1_1772(.clk(clk),.reset(reset),.i1(intermediate_reg_0[55]),.i2(intermediate_reg_0[54]),.o(intermediate_reg_1[27]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1773(.clk(clk),.reset(reset),.i1(intermediate_reg_0[53]),.i2(intermediate_reg_0[52]),.o(intermediate_reg_1[26])); 
mux_module mux_module_inst_1_1774(.clk(clk),.reset(reset),.i1(intermediate_reg_0[51]),.i2(intermediate_reg_0[50]),.o(intermediate_reg_1[25]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1775(.clk(clk),.reset(reset),.i1(intermediate_reg_0[49]),.i2(intermediate_reg_0[48]),.o(intermediate_reg_1[24])); 
fsm fsm_inst_1_1776(.clk(clk),.reset(reset),.i1(intermediate_reg_0[47]),.i2(intermediate_reg_0[46]),.o(intermediate_reg_1[23])); 
fsm fsm_inst_1_1777(.clk(clk),.reset(reset),.i1(intermediate_reg_0[45]),.i2(intermediate_reg_0[44]),.o(intermediate_reg_1[22])); 
fsm fsm_inst_1_1778(.clk(clk),.reset(reset),.i1(intermediate_reg_0[43]),.i2(intermediate_reg_0[42]),.o(intermediate_reg_1[21])); 
mux_module mux_module_inst_1_1779(.clk(clk),.reset(reset),.i1(intermediate_reg_0[41]),.i2(intermediate_reg_0[40]),.o(intermediate_reg_1[20]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1780(.clk(clk),.reset(reset),.i1(intermediate_reg_0[39]),.i2(intermediate_reg_0[38]),.o(intermediate_reg_1[19])); 
mux_module mux_module_inst_1_1781(.clk(clk),.reset(reset),.i1(intermediate_reg_0[37]),.i2(intermediate_reg_0[36]),.o(intermediate_reg_1[18]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1782(.clk(clk),.reset(reset),.i1(intermediate_reg_0[35]),.i2(intermediate_reg_0[34]),.o(intermediate_reg_1[17]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1783(.clk(clk),.reset(reset),.i1(intermediate_reg_0[33]),.i2(intermediate_reg_0[32]),.o(intermediate_reg_1[16]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1784(.clk(clk),.reset(reset),.i1(intermediate_reg_0[31]),.i2(intermediate_reg_0[30]),.o(intermediate_reg_1[15])); 
mux_module mux_module_inst_1_1785(.clk(clk),.reset(reset),.i1(intermediate_reg_0[29]),.i2(intermediate_reg_0[28]),.o(intermediate_reg_1[14]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1786(.clk(clk),.reset(reset),.i1(intermediate_reg_0[27]),.i2(intermediate_reg_0[26]),.o(intermediate_reg_1[13]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1787(.clk(clk),.reset(reset),.i1(intermediate_reg_0[25]),.i2(intermediate_reg_0[24]),.o(intermediate_reg_1[12]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1788(.clk(clk),.reset(reset),.i1(intermediate_reg_0[23]),.i2(intermediate_reg_0[22]),.o(intermediate_reg_1[11]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1789(.clk(clk),.reset(reset),.i1(intermediate_reg_0[21]),.i2(intermediate_reg_0[20]),.o(intermediate_reg_1[10]),.sel(intermediate_reg_0[0])); 
mux_module mux_module_inst_1_1790(.clk(clk),.reset(reset),.i1(intermediate_reg_0[19]),.i2(intermediate_reg_0[18]),.o(intermediate_reg_1[9]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1791(.clk(clk),.reset(reset),.i1(intermediate_reg_0[17]),.i2(intermediate_reg_0[16]),.o(intermediate_reg_1[8])); 
fsm fsm_inst_1_1792(.clk(clk),.reset(reset),.i1(intermediate_reg_0[15]),.i2(intermediate_reg_0[14]),.o(intermediate_reg_1[7])); 
fsm fsm_inst_1_1793(.clk(clk),.reset(reset),.i1(intermediate_reg_0[13]),.i2(intermediate_reg_0[12]),.o(intermediate_reg_1[6])); 
fsm fsm_inst_1_1794(.clk(clk),.reset(reset),.i1(intermediate_reg_0[11]),.i2(intermediate_reg_0[10]),.o(intermediate_reg_1[5])); 
fsm fsm_inst_1_1795(.clk(clk),.reset(reset),.i1(intermediate_reg_0[9]),.i2(intermediate_reg_0[8]),.o(intermediate_reg_1[4])); 
fsm fsm_inst_1_1796(.clk(clk),.reset(reset),.i1(intermediate_reg_0[7]),.i2(intermediate_reg_0[6]),.o(intermediate_reg_1[3])); 
mux_module mux_module_inst_1_1797(.clk(clk),.reset(reset),.i1(intermediate_reg_0[5]),.i2(intermediate_reg_0[4]),.o(intermediate_reg_1[2]),.sel(intermediate_reg_0[0])); 
fsm fsm_inst_1_1798(.clk(clk),.reset(reset),.i1(intermediate_reg_0[3]),.i2(intermediate_reg_0[2]),.o(intermediate_reg_1[1])); 
mux_module mux_module_inst_1_1799(.clk(clk),.reset(reset),.i1(intermediate_reg_0[1]),.i2(intermediate_reg_0[0]),.o(intermediate_reg_1[0]),.sel(intermediate_reg_0[0])); 
reg [899:0]intermediate_reg_2; 
 
mux_module mux_module_inst_2_0(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1799]),.i2(intermediate_reg_1[1798]),.o(intermediate_reg_2[899]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_1(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1797]),.i2(intermediate_reg_1[1796]),.o(intermediate_reg_2[898]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_2(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1795]),.i2(intermediate_reg_1[1794]),.o(intermediate_reg_2[897]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_3(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1793]),.i2(intermediate_reg_1[1792]),.o(intermediate_reg_2[896]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_4(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1791]),.i2(intermediate_reg_1[1790]),.o(intermediate_reg_2[895])); 
mux_module mux_module_inst_2_5(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1789]),.i2(intermediate_reg_1[1788]),.o(intermediate_reg_2[894]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_6(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1787]),.i2(intermediate_reg_1[1786]),.o(intermediate_reg_2[893]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_7(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1785]),.i2(intermediate_reg_1[1784]),.o(intermediate_reg_2[892]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_8(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1783]),.i2(intermediate_reg_1[1782]),.o(intermediate_reg_2[891]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_9(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1781]),.i2(intermediate_reg_1[1780]),.o(intermediate_reg_2[890]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_10(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1779]),.i2(intermediate_reg_1[1778]),.o(intermediate_reg_2[889])); 
mux_module mux_module_inst_2_11(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1777]),.i2(intermediate_reg_1[1776]),.o(intermediate_reg_2[888]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_12(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1775]),.i2(intermediate_reg_1[1774]),.o(intermediate_reg_2[887])); 
mux_module mux_module_inst_2_13(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1773]),.i2(intermediate_reg_1[1772]),.o(intermediate_reg_2[886]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_14(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1771]),.i2(intermediate_reg_1[1770]),.o(intermediate_reg_2[885]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_15(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1769]),.i2(intermediate_reg_1[1768]),.o(intermediate_reg_2[884]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_16(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1767]),.i2(intermediate_reg_1[1766]),.o(intermediate_reg_2[883]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_17(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1765]),.i2(intermediate_reg_1[1764]),.o(intermediate_reg_2[882]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_18(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1763]),.i2(intermediate_reg_1[1762]),.o(intermediate_reg_2[881]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_19(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1761]),.i2(intermediate_reg_1[1760]),.o(intermediate_reg_2[880]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_20(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1759]),.i2(intermediate_reg_1[1758]),.o(intermediate_reg_2[879])); 
fsm fsm_inst_2_21(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1757]),.i2(intermediate_reg_1[1756]),.o(intermediate_reg_2[878])); 
fsm fsm_inst_2_22(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1755]),.i2(intermediate_reg_1[1754]),.o(intermediate_reg_2[877])); 
fsm fsm_inst_2_23(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1753]),.i2(intermediate_reg_1[1752]),.o(intermediate_reg_2[876])); 
fsm fsm_inst_2_24(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1751]),.i2(intermediate_reg_1[1750]),.o(intermediate_reg_2[875])); 
fsm fsm_inst_2_25(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1749]),.i2(intermediate_reg_1[1748]),.o(intermediate_reg_2[874])); 
mux_module mux_module_inst_2_26(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1747]),.i2(intermediate_reg_1[1746]),.o(intermediate_reg_2[873]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_27(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1745]),.i2(intermediate_reg_1[1744]),.o(intermediate_reg_2[872])); 
mux_module mux_module_inst_2_28(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1743]),.i2(intermediate_reg_1[1742]),.o(intermediate_reg_2[871]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_29(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1741]),.i2(intermediate_reg_1[1740]),.o(intermediate_reg_2[870]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_30(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1739]),.i2(intermediate_reg_1[1738]),.o(intermediate_reg_2[869])); 
fsm fsm_inst_2_31(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1737]),.i2(intermediate_reg_1[1736]),.o(intermediate_reg_2[868])); 
fsm fsm_inst_2_32(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1735]),.i2(intermediate_reg_1[1734]),.o(intermediate_reg_2[867])); 
fsm fsm_inst_2_33(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1733]),.i2(intermediate_reg_1[1732]),.o(intermediate_reg_2[866])); 
fsm fsm_inst_2_34(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1731]),.i2(intermediate_reg_1[1730]),.o(intermediate_reg_2[865])); 
mux_module mux_module_inst_2_35(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1729]),.i2(intermediate_reg_1[1728]),.o(intermediate_reg_2[864]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_36(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1727]),.i2(intermediate_reg_1[1726]),.o(intermediate_reg_2[863])); 
mux_module mux_module_inst_2_37(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1725]),.i2(intermediate_reg_1[1724]),.o(intermediate_reg_2[862]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_38(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1723]),.i2(intermediate_reg_1[1722]),.o(intermediate_reg_2[861]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_39(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1721]),.i2(intermediate_reg_1[1720]),.o(intermediate_reg_2[860]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_40(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1719]),.i2(intermediate_reg_1[1718]),.o(intermediate_reg_2[859])); 
mux_module mux_module_inst_2_41(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1717]),.i2(intermediate_reg_1[1716]),.o(intermediate_reg_2[858]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_42(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1715]),.i2(intermediate_reg_1[1714]),.o(intermediate_reg_2[857]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_43(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1713]),.i2(intermediate_reg_1[1712]),.o(intermediate_reg_2[856])); 
mux_module mux_module_inst_2_44(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1711]),.i2(intermediate_reg_1[1710]),.o(intermediate_reg_2[855]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_45(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1709]),.i2(intermediate_reg_1[1708]),.o(intermediate_reg_2[854])); 
fsm fsm_inst_2_46(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1707]),.i2(intermediate_reg_1[1706]),.o(intermediate_reg_2[853])); 
mux_module mux_module_inst_2_47(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1705]),.i2(intermediate_reg_1[1704]),.o(intermediate_reg_2[852]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_48(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1703]),.i2(intermediate_reg_1[1702]),.o(intermediate_reg_2[851])); 
mux_module mux_module_inst_2_49(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1701]),.i2(intermediate_reg_1[1700]),.o(intermediate_reg_2[850]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_50(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1699]),.i2(intermediate_reg_1[1698]),.o(intermediate_reg_2[849]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_51(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1697]),.i2(intermediate_reg_1[1696]),.o(intermediate_reg_2[848]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_52(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1695]),.i2(intermediate_reg_1[1694]),.o(intermediate_reg_2[847])); 
mux_module mux_module_inst_2_53(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1693]),.i2(intermediate_reg_1[1692]),.o(intermediate_reg_2[846]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_54(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1691]),.i2(intermediate_reg_1[1690]),.o(intermediate_reg_2[845]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_55(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1689]),.i2(intermediate_reg_1[1688]),.o(intermediate_reg_2[844]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_56(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1687]),.i2(intermediate_reg_1[1686]),.o(intermediate_reg_2[843])); 
mux_module mux_module_inst_2_57(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1685]),.i2(intermediate_reg_1[1684]),.o(intermediate_reg_2[842]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_58(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1683]),.i2(intermediate_reg_1[1682]),.o(intermediate_reg_2[841])); 
mux_module mux_module_inst_2_59(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1681]),.i2(intermediate_reg_1[1680]),.o(intermediate_reg_2[840]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_60(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1679]),.i2(intermediate_reg_1[1678]),.o(intermediate_reg_2[839]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_61(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1677]),.i2(intermediate_reg_1[1676]),.o(intermediate_reg_2[838])); 
fsm fsm_inst_2_62(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1675]),.i2(intermediate_reg_1[1674]),.o(intermediate_reg_2[837])); 
fsm fsm_inst_2_63(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1673]),.i2(intermediate_reg_1[1672]),.o(intermediate_reg_2[836])); 
fsm fsm_inst_2_64(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1671]),.i2(intermediate_reg_1[1670]),.o(intermediate_reg_2[835])); 
fsm fsm_inst_2_65(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1669]),.i2(intermediate_reg_1[1668]),.o(intermediate_reg_2[834])); 
mux_module mux_module_inst_2_66(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1667]),.i2(intermediate_reg_1[1666]),.o(intermediate_reg_2[833]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_67(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1665]),.i2(intermediate_reg_1[1664]),.o(intermediate_reg_2[832]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_68(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1663]),.i2(intermediate_reg_1[1662]),.o(intermediate_reg_2[831]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_69(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1661]),.i2(intermediate_reg_1[1660]),.o(intermediate_reg_2[830])); 
fsm fsm_inst_2_70(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1659]),.i2(intermediate_reg_1[1658]),.o(intermediate_reg_2[829])); 
mux_module mux_module_inst_2_71(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1657]),.i2(intermediate_reg_1[1656]),.o(intermediate_reg_2[828]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_72(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1655]),.i2(intermediate_reg_1[1654]),.o(intermediate_reg_2[827])); 
fsm fsm_inst_2_73(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1653]),.i2(intermediate_reg_1[1652]),.o(intermediate_reg_2[826])); 
fsm fsm_inst_2_74(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1651]),.i2(intermediate_reg_1[1650]),.o(intermediate_reg_2[825])); 
fsm fsm_inst_2_75(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1649]),.i2(intermediate_reg_1[1648]),.o(intermediate_reg_2[824])); 
mux_module mux_module_inst_2_76(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1647]),.i2(intermediate_reg_1[1646]),.o(intermediate_reg_2[823]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_77(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1645]),.i2(intermediate_reg_1[1644]),.o(intermediate_reg_2[822]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_78(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1643]),.i2(intermediate_reg_1[1642]),.o(intermediate_reg_2[821])); 
fsm fsm_inst_2_79(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1641]),.i2(intermediate_reg_1[1640]),.o(intermediate_reg_2[820])); 
fsm fsm_inst_2_80(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1639]),.i2(intermediate_reg_1[1638]),.o(intermediate_reg_2[819])); 
mux_module mux_module_inst_2_81(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1637]),.i2(intermediate_reg_1[1636]),.o(intermediate_reg_2[818]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_82(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1635]),.i2(intermediate_reg_1[1634]),.o(intermediate_reg_2[817]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_83(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1633]),.i2(intermediate_reg_1[1632]),.o(intermediate_reg_2[816])); 
fsm fsm_inst_2_84(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1631]),.i2(intermediate_reg_1[1630]),.o(intermediate_reg_2[815])); 
fsm fsm_inst_2_85(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1629]),.i2(intermediate_reg_1[1628]),.o(intermediate_reg_2[814])); 
mux_module mux_module_inst_2_86(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1627]),.i2(intermediate_reg_1[1626]),.o(intermediate_reg_2[813]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_87(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1625]),.i2(intermediate_reg_1[1624]),.o(intermediate_reg_2[812])); 
mux_module mux_module_inst_2_88(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1623]),.i2(intermediate_reg_1[1622]),.o(intermediate_reg_2[811]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_89(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1621]),.i2(intermediate_reg_1[1620]),.o(intermediate_reg_2[810])); 
mux_module mux_module_inst_2_90(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1619]),.i2(intermediate_reg_1[1618]),.o(intermediate_reg_2[809]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_91(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1617]),.i2(intermediate_reg_1[1616]),.o(intermediate_reg_2[808]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_92(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1615]),.i2(intermediate_reg_1[1614]),.o(intermediate_reg_2[807])); 
fsm fsm_inst_2_93(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1613]),.i2(intermediate_reg_1[1612]),.o(intermediate_reg_2[806])); 
fsm fsm_inst_2_94(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1611]),.i2(intermediate_reg_1[1610]),.o(intermediate_reg_2[805])); 
mux_module mux_module_inst_2_95(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1609]),.i2(intermediate_reg_1[1608]),.o(intermediate_reg_2[804]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_96(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1607]),.i2(intermediate_reg_1[1606]),.o(intermediate_reg_2[803]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_97(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1605]),.i2(intermediate_reg_1[1604]),.o(intermediate_reg_2[802])); 
mux_module mux_module_inst_2_98(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1603]),.i2(intermediate_reg_1[1602]),.o(intermediate_reg_2[801]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_99(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1601]),.i2(intermediate_reg_1[1600]),.o(intermediate_reg_2[800])); 
fsm fsm_inst_2_100(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1599]),.i2(intermediate_reg_1[1598]),.o(intermediate_reg_2[799])); 
fsm fsm_inst_2_101(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1597]),.i2(intermediate_reg_1[1596]),.o(intermediate_reg_2[798])); 
mux_module mux_module_inst_2_102(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1595]),.i2(intermediate_reg_1[1594]),.o(intermediate_reg_2[797]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_103(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1593]),.i2(intermediate_reg_1[1592]),.o(intermediate_reg_2[796]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_104(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1591]),.i2(intermediate_reg_1[1590]),.o(intermediate_reg_2[795]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_105(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1589]),.i2(intermediate_reg_1[1588]),.o(intermediate_reg_2[794])); 
fsm fsm_inst_2_106(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1587]),.i2(intermediate_reg_1[1586]),.o(intermediate_reg_2[793])); 
fsm fsm_inst_2_107(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1585]),.i2(intermediate_reg_1[1584]),.o(intermediate_reg_2[792])); 
mux_module mux_module_inst_2_108(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1583]),.i2(intermediate_reg_1[1582]),.o(intermediate_reg_2[791]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_109(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1581]),.i2(intermediate_reg_1[1580]),.o(intermediate_reg_2[790])); 
fsm fsm_inst_2_110(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1579]),.i2(intermediate_reg_1[1578]),.o(intermediate_reg_2[789])); 
mux_module mux_module_inst_2_111(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1577]),.i2(intermediate_reg_1[1576]),.o(intermediate_reg_2[788]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_112(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1575]),.i2(intermediate_reg_1[1574]),.o(intermediate_reg_2[787]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_113(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1573]),.i2(intermediate_reg_1[1572]),.o(intermediate_reg_2[786]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_114(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1571]),.i2(intermediate_reg_1[1570]),.o(intermediate_reg_2[785])); 
fsm fsm_inst_2_115(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1569]),.i2(intermediate_reg_1[1568]),.o(intermediate_reg_2[784])); 
mux_module mux_module_inst_2_116(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1567]),.i2(intermediate_reg_1[1566]),.o(intermediate_reg_2[783]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_117(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1565]),.i2(intermediate_reg_1[1564]),.o(intermediate_reg_2[782])); 
mux_module mux_module_inst_2_118(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1563]),.i2(intermediate_reg_1[1562]),.o(intermediate_reg_2[781]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_119(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1561]),.i2(intermediate_reg_1[1560]),.o(intermediate_reg_2[780]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_120(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1559]),.i2(intermediate_reg_1[1558]),.o(intermediate_reg_2[779]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_121(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1557]),.i2(intermediate_reg_1[1556]),.o(intermediate_reg_2[778])); 
mux_module mux_module_inst_2_122(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1555]),.i2(intermediate_reg_1[1554]),.o(intermediate_reg_2[777]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_123(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1553]),.i2(intermediate_reg_1[1552]),.o(intermediate_reg_2[776])); 
fsm fsm_inst_2_124(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1551]),.i2(intermediate_reg_1[1550]),.o(intermediate_reg_2[775])); 
fsm fsm_inst_2_125(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1549]),.i2(intermediate_reg_1[1548]),.o(intermediate_reg_2[774])); 
mux_module mux_module_inst_2_126(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1547]),.i2(intermediate_reg_1[1546]),.o(intermediate_reg_2[773]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_127(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1545]),.i2(intermediate_reg_1[1544]),.o(intermediate_reg_2[772]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_128(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1543]),.i2(intermediate_reg_1[1542]),.o(intermediate_reg_2[771])); 
fsm fsm_inst_2_129(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1541]),.i2(intermediate_reg_1[1540]),.o(intermediate_reg_2[770])); 
fsm fsm_inst_2_130(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1539]),.i2(intermediate_reg_1[1538]),.o(intermediate_reg_2[769])); 
fsm fsm_inst_2_131(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1537]),.i2(intermediate_reg_1[1536]),.o(intermediate_reg_2[768])); 
mux_module mux_module_inst_2_132(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1535]),.i2(intermediate_reg_1[1534]),.o(intermediate_reg_2[767]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_133(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1533]),.i2(intermediate_reg_1[1532]),.o(intermediate_reg_2[766]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_134(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1531]),.i2(intermediate_reg_1[1530]),.o(intermediate_reg_2[765]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_135(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1529]),.i2(intermediate_reg_1[1528]),.o(intermediate_reg_2[764]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_136(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1527]),.i2(intermediate_reg_1[1526]),.o(intermediate_reg_2[763]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_137(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1525]),.i2(intermediate_reg_1[1524]),.o(intermediate_reg_2[762]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_138(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1523]),.i2(intermediate_reg_1[1522]),.o(intermediate_reg_2[761])); 
fsm fsm_inst_2_139(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1521]),.i2(intermediate_reg_1[1520]),.o(intermediate_reg_2[760])); 
mux_module mux_module_inst_2_140(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1519]),.i2(intermediate_reg_1[1518]),.o(intermediate_reg_2[759]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_141(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1517]),.i2(intermediate_reg_1[1516]),.o(intermediate_reg_2[758])); 
fsm fsm_inst_2_142(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1515]),.i2(intermediate_reg_1[1514]),.o(intermediate_reg_2[757])); 
fsm fsm_inst_2_143(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1513]),.i2(intermediate_reg_1[1512]),.o(intermediate_reg_2[756])); 
mux_module mux_module_inst_2_144(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1511]),.i2(intermediate_reg_1[1510]),.o(intermediate_reg_2[755]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_145(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1509]),.i2(intermediate_reg_1[1508]),.o(intermediate_reg_2[754])); 
mux_module mux_module_inst_2_146(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1507]),.i2(intermediate_reg_1[1506]),.o(intermediate_reg_2[753]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_147(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1505]),.i2(intermediate_reg_1[1504]),.o(intermediate_reg_2[752]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_148(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1503]),.i2(intermediate_reg_1[1502]),.o(intermediate_reg_2[751])); 
mux_module mux_module_inst_2_149(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1501]),.i2(intermediate_reg_1[1500]),.o(intermediate_reg_2[750]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_150(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1499]),.i2(intermediate_reg_1[1498]),.o(intermediate_reg_2[749]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_151(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1497]),.i2(intermediate_reg_1[1496]),.o(intermediate_reg_2[748]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_152(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1495]),.i2(intermediate_reg_1[1494]),.o(intermediate_reg_2[747]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_153(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1493]),.i2(intermediate_reg_1[1492]),.o(intermediate_reg_2[746])); 
fsm fsm_inst_2_154(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1491]),.i2(intermediate_reg_1[1490]),.o(intermediate_reg_2[745])); 
fsm fsm_inst_2_155(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1489]),.i2(intermediate_reg_1[1488]),.o(intermediate_reg_2[744])); 
fsm fsm_inst_2_156(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1487]),.i2(intermediate_reg_1[1486]),.o(intermediate_reg_2[743])); 
fsm fsm_inst_2_157(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1485]),.i2(intermediate_reg_1[1484]),.o(intermediate_reg_2[742])); 
fsm fsm_inst_2_158(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1483]),.i2(intermediate_reg_1[1482]),.o(intermediate_reg_2[741])); 
mux_module mux_module_inst_2_159(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1481]),.i2(intermediate_reg_1[1480]),.o(intermediate_reg_2[740]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_160(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1479]),.i2(intermediate_reg_1[1478]),.o(intermediate_reg_2[739]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_161(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1477]),.i2(intermediate_reg_1[1476]),.o(intermediate_reg_2[738])); 
fsm fsm_inst_2_162(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1475]),.i2(intermediate_reg_1[1474]),.o(intermediate_reg_2[737])); 
fsm fsm_inst_2_163(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1473]),.i2(intermediate_reg_1[1472]),.o(intermediate_reg_2[736])); 
mux_module mux_module_inst_2_164(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1471]),.i2(intermediate_reg_1[1470]),.o(intermediate_reg_2[735]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_165(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1469]),.i2(intermediate_reg_1[1468]),.o(intermediate_reg_2[734])); 
mux_module mux_module_inst_2_166(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1467]),.i2(intermediate_reg_1[1466]),.o(intermediate_reg_2[733]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_167(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1465]),.i2(intermediate_reg_1[1464]),.o(intermediate_reg_2[732])); 
mux_module mux_module_inst_2_168(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1463]),.i2(intermediate_reg_1[1462]),.o(intermediate_reg_2[731]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_169(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1461]),.i2(intermediate_reg_1[1460]),.o(intermediate_reg_2[730])); 
mux_module mux_module_inst_2_170(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1459]),.i2(intermediate_reg_1[1458]),.o(intermediate_reg_2[729]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_171(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1457]),.i2(intermediate_reg_1[1456]),.o(intermediate_reg_2[728]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_172(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1455]),.i2(intermediate_reg_1[1454]),.o(intermediate_reg_2[727]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_173(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1453]),.i2(intermediate_reg_1[1452]),.o(intermediate_reg_2[726])); 
mux_module mux_module_inst_2_174(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1451]),.i2(intermediate_reg_1[1450]),.o(intermediate_reg_2[725]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_175(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1449]),.i2(intermediate_reg_1[1448]),.o(intermediate_reg_2[724]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_176(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1447]),.i2(intermediate_reg_1[1446]),.o(intermediate_reg_2[723])); 
fsm fsm_inst_2_177(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1445]),.i2(intermediate_reg_1[1444]),.o(intermediate_reg_2[722])); 
fsm fsm_inst_2_178(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1443]),.i2(intermediate_reg_1[1442]),.o(intermediate_reg_2[721])); 
fsm fsm_inst_2_179(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1441]),.i2(intermediate_reg_1[1440]),.o(intermediate_reg_2[720])); 
mux_module mux_module_inst_2_180(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1439]),.i2(intermediate_reg_1[1438]),.o(intermediate_reg_2[719]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_181(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1437]),.i2(intermediate_reg_1[1436]),.o(intermediate_reg_2[718]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_182(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1435]),.i2(intermediate_reg_1[1434]),.o(intermediate_reg_2[717]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_183(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1433]),.i2(intermediate_reg_1[1432]),.o(intermediate_reg_2[716])); 
fsm fsm_inst_2_184(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1431]),.i2(intermediate_reg_1[1430]),.o(intermediate_reg_2[715])); 
mux_module mux_module_inst_2_185(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1429]),.i2(intermediate_reg_1[1428]),.o(intermediate_reg_2[714]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_186(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1427]),.i2(intermediate_reg_1[1426]),.o(intermediate_reg_2[713])); 
mux_module mux_module_inst_2_187(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1425]),.i2(intermediate_reg_1[1424]),.o(intermediate_reg_2[712]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_188(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1423]),.i2(intermediate_reg_1[1422]),.o(intermediate_reg_2[711]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_189(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1421]),.i2(intermediate_reg_1[1420]),.o(intermediate_reg_2[710])); 
fsm fsm_inst_2_190(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1419]),.i2(intermediate_reg_1[1418]),.o(intermediate_reg_2[709])); 
fsm fsm_inst_2_191(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1417]),.i2(intermediate_reg_1[1416]),.o(intermediate_reg_2[708])); 
mux_module mux_module_inst_2_192(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1415]),.i2(intermediate_reg_1[1414]),.o(intermediate_reg_2[707]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_193(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1413]),.i2(intermediate_reg_1[1412]),.o(intermediate_reg_2[706])); 
fsm fsm_inst_2_194(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1411]),.i2(intermediate_reg_1[1410]),.o(intermediate_reg_2[705])); 
fsm fsm_inst_2_195(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1409]),.i2(intermediate_reg_1[1408]),.o(intermediate_reg_2[704])); 
mux_module mux_module_inst_2_196(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1407]),.i2(intermediate_reg_1[1406]),.o(intermediate_reg_2[703]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_197(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1405]),.i2(intermediate_reg_1[1404]),.o(intermediate_reg_2[702])); 
mux_module mux_module_inst_2_198(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1403]),.i2(intermediate_reg_1[1402]),.o(intermediate_reg_2[701]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_199(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1401]),.i2(intermediate_reg_1[1400]),.o(intermediate_reg_2[700])); 
mux_module mux_module_inst_2_200(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1399]),.i2(intermediate_reg_1[1398]),.o(intermediate_reg_2[699]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_201(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1397]),.i2(intermediate_reg_1[1396]),.o(intermediate_reg_2[698]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_202(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1395]),.i2(intermediate_reg_1[1394]),.o(intermediate_reg_2[697])); 
mux_module mux_module_inst_2_203(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1393]),.i2(intermediate_reg_1[1392]),.o(intermediate_reg_2[696]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_204(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1391]),.i2(intermediate_reg_1[1390]),.o(intermediate_reg_2[695]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_205(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1389]),.i2(intermediate_reg_1[1388]),.o(intermediate_reg_2[694]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_206(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1387]),.i2(intermediate_reg_1[1386]),.o(intermediate_reg_2[693])); 
mux_module mux_module_inst_2_207(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1385]),.i2(intermediate_reg_1[1384]),.o(intermediate_reg_2[692]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_208(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1383]),.i2(intermediate_reg_1[1382]),.o(intermediate_reg_2[691])); 
fsm fsm_inst_2_209(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1381]),.i2(intermediate_reg_1[1380]),.o(intermediate_reg_2[690])); 
mux_module mux_module_inst_2_210(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1379]),.i2(intermediate_reg_1[1378]),.o(intermediate_reg_2[689]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_211(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1377]),.i2(intermediate_reg_1[1376]),.o(intermediate_reg_2[688]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_212(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1375]),.i2(intermediate_reg_1[1374]),.o(intermediate_reg_2[687])); 
mux_module mux_module_inst_2_213(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1373]),.i2(intermediate_reg_1[1372]),.o(intermediate_reg_2[686]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_214(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1371]),.i2(intermediate_reg_1[1370]),.o(intermediate_reg_2[685]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_215(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1369]),.i2(intermediate_reg_1[1368]),.o(intermediate_reg_2[684])); 
fsm fsm_inst_2_216(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1367]),.i2(intermediate_reg_1[1366]),.o(intermediate_reg_2[683])); 
mux_module mux_module_inst_2_217(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1365]),.i2(intermediate_reg_1[1364]),.o(intermediate_reg_2[682]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_218(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1363]),.i2(intermediate_reg_1[1362]),.o(intermediate_reg_2[681]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_219(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1361]),.i2(intermediate_reg_1[1360]),.o(intermediate_reg_2[680])); 
fsm fsm_inst_2_220(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1359]),.i2(intermediate_reg_1[1358]),.o(intermediate_reg_2[679])); 
fsm fsm_inst_2_221(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1357]),.i2(intermediate_reg_1[1356]),.o(intermediate_reg_2[678])); 
fsm fsm_inst_2_222(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1355]),.i2(intermediate_reg_1[1354]),.o(intermediate_reg_2[677])); 
fsm fsm_inst_2_223(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1353]),.i2(intermediate_reg_1[1352]),.o(intermediate_reg_2[676])); 
fsm fsm_inst_2_224(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1351]),.i2(intermediate_reg_1[1350]),.o(intermediate_reg_2[675])); 
mux_module mux_module_inst_2_225(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1349]),.i2(intermediate_reg_1[1348]),.o(intermediate_reg_2[674]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_226(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1347]),.i2(intermediate_reg_1[1346]),.o(intermediate_reg_2[673]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_227(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1345]),.i2(intermediate_reg_1[1344]),.o(intermediate_reg_2[672])); 
mux_module mux_module_inst_2_228(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1343]),.i2(intermediate_reg_1[1342]),.o(intermediate_reg_2[671]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_229(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1341]),.i2(intermediate_reg_1[1340]),.o(intermediate_reg_2[670])); 
fsm fsm_inst_2_230(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1339]),.i2(intermediate_reg_1[1338]),.o(intermediate_reg_2[669])); 
mux_module mux_module_inst_2_231(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1337]),.i2(intermediate_reg_1[1336]),.o(intermediate_reg_2[668]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_232(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1335]),.i2(intermediate_reg_1[1334]),.o(intermediate_reg_2[667])); 
fsm fsm_inst_2_233(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1333]),.i2(intermediate_reg_1[1332]),.o(intermediate_reg_2[666])); 
fsm fsm_inst_2_234(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1331]),.i2(intermediate_reg_1[1330]),.o(intermediate_reg_2[665])); 
fsm fsm_inst_2_235(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1329]),.i2(intermediate_reg_1[1328]),.o(intermediate_reg_2[664])); 
mux_module mux_module_inst_2_236(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1327]),.i2(intermediate_reg_1[1326]),.o(intermediate_reg_2[663]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_237(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1325]),.i2(intermediate_reg_1[1324]),.o(intermediate_reg_2[662]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_238(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1323]),.i2(intermediate_reg_1[1322]),.o(intermediate_reg_2[661]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_239(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1321]),.i2(intermediate_reg_1[1320]),.o(intermediate_reg_2[660])); 
fsm fsm_inst_2_240(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1319]),.i2(intermediate_reg_1[1318]),.o(intermediate_reg_2[659])); 
fsm fsm_inst_2_241(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1317]),.i2(intermediate_reg_1[1316]),.o(intermediate_reg_2[658])); 
fsm fsm_inst_2_242(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1315]),.i2(intermediate_reg_1[1314]),.o(intermediate_reg_2[657])); 
mux_module mux_module_inst_2_243(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1313]),.i2(intermediate_reg_1[1312]),.o(intermediate_reg_2[656]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_244(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1311]),.i2(intermediate_reg_1[1310]),.o(intermediate_reg_2[655]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_245(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1309]),.i2(intermediate_reg_1[1308]),.o(intermediate_reg_2[654])); 
fsm fsm_inst_2_246(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1307]),.i2(intermediate_reg_1[1306]),.o(intermediate_reg_2[653])); 
fsm fsm_inst_2_247(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1305]),.i2(intermediate_reg_1[1304]),.o(intermediate_reg_2[652])); 
fsm fsm_inst_2_248(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1303]),.i2(intermediate_reg_1[1302]),.o(intermediate_reg_2[651])); 
fsm fsm_inst_2_249(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1301]),.i2(intermediate_reg_1[1300]),.o(intermediate_reg_2[650])); 
mux_module mux_module_inst_2_250(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1299]),.i2(intermediate_reg_1[1298]),.o(intermediate_reg_2[649]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_251(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1297]),.i2(intermediate_reg_1[1296]),.o(intermediate_reg_2[648])); 
mux_module mux_module_inst_2_252(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1295]),.i2(intermediate_reg_1[1294]),.o(intermediate_reg_2[647]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_253(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1293]),.i2(intermediate_reg_1[1292]),.o(intermediate_reg_2[646]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_254(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1291]),.i2(intermediate_reg_1[1290]),.o(intermediate_reg_2[645])); 
fsm fsm_inst_2_255(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1289]),.i2(intermediate_reg_1[1288]),.o(intermediate_reg_2[644])); 
fsm fsm_inst_2_256(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1287]),.i2(intermediate_reg_1[1286]),.o(intermediate_reg_2[643])); 
mux_module mux_module_inst_2_257(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1285]),.i2(intermediate_reg_1[1284]),.o(intermediate_reg_2[642]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_258(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1283]),.i2(intermediate_reg_1[1282]),.o(intermediate_reg_2[641]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_259(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1281]),.i2(intermediate_reg_1[1280]),.o(intermediate_reg_2[640]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_260(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1279]),.i2(intermediate_reg_1[1278]),.o(intermediate_reg_2[639]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_261(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1277]),.i2(intermediate_reg_1[1276]),.o(intermediate_reg_2[638])); 
fsm fsm_inst_2_262(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1275]),.i2(intermediate_reg_1[1274]),.o(intermediate_reg_2[637])); 
mux_module mux_module_inst_2_263(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1273]),.i2(intermediate_reg_1[1272]),.o(intermediate_reg_2[636]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_264(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1271]),.i2(intermediate_reg_1[1270]),.o(intermediate_reg_2[635])); 
mux_module mux_module_inst_2_265(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1269]),.i2(intermediate_reg_1[1268]),.o(intermediate_reg_2[634]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_266(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1267]),.i2(intermediate_reg_1[1266]),.o(intermediate_reg_2[633])); 
fsm fsm_inst_2_267(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1265]),.i2(intermediate_reg_1[1264]),.o(intermediate_reg_2[632])); 
mux_module mux_module_inst_2_268(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1263]),.i2(intermediate_reg_1[1262]),.o(intermediate_reg_2[631]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_269(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1261]),.i2(intermediate_reg_1[1260]),.o(intermediate_reg_2[630])); 
fsm fsm_inst_2_270(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1259]),.i2(intermediate_reg_1[1258]),.o(intermediate_reg_2[629])); 
fsm fsm_inst_2_271(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1257]),.i2(intermediate_reg_1[1256]),.o(intermediate_reg_2[628])); 
mux_module mux_module_inst_2_272(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1255]),.i2(intermediate_reg_1[1254]),.o(intermediate_reg_2[627]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_273(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1253]),.i2(intermediate_reg_1[1252]),.o(intermediate_reg_2[626]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_274(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1251]),.i2(intermediate_reg_1[1250]),.o(intermediate_reg_2[625])); 
mux_module mux_module_inst_2_275(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1249]),.i2(intermediate_reg_1[1248]),.o(intermediate_reg_2[624]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_276(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1247]),.i2(intermediate_reg_1[1246]),.o(intermediate_reg_2[623]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_277(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1245]),.i2(intermediate_reg_1[1244]),.o(intermediate_reg_2[622])); 
fsm fsm_inst_2_278(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1243]),.i2(intermediate_reg_1[1242]),.o(intermediate_reg_2[621])); 
fsm fsm_inst_2_279(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1241]),.i2(intermediate_reg_1[1240]),.o(intermediate_reg_2[620])); 
fsm fsm_inst_2_280(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1239]),.i2(intermediate_reg_1[1238]),.o(intermediate_reg_2[619])); 
mux_module mux_module_inst_2_281(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1237]),.i2(intermediate_reg_1[1236]),.o(intermediate_reg_2[618]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_282(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1235]),.i2(intermediate_reg_1[1234]),.o(intermediate_reg_2[617]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_283(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1233]),.i2(intermediate_reg_1[1232]),.o(intermediate_reg_2[616]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_284(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1231]),.i2(intermediate_reg_1[1230]),.o(intermediate_reg_2[615]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_285(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1229]),.i2(intermediate_reg_1[1228]),.o(intermediate_reg_2[614]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_286(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1227]),.i2(intermediate_reg_1[1226]),.o(intermediate_reg_2[613])); 
fsm fsm_inst_2_287(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1225]),.i2(intermediate_reg_1[1224]),.o(intermediate_reg_2[612])); 
fsm fsm_inst_2_288(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1223]),.i2(intermediate_reg_1[1222]),.o(intermediate_reg_2[611])); 
mux_module mux_module_inst_2_289(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1221]),.i2(intermediate_reg_1[1220]),.o(intermediate_reg_2[610]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_290(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1219]),.i2(intermediate_reg_1[1218]),.o(intermediate_reg_2[609])); 
fsm fsm_inst_2_291(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1217]),.i2(intermediate_reg_1[1216]),.o(intermediate_reg_2[608])); 
fsm fsm_inst_2_292(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1215]),.i2(intermediate_reg_1[1214]),.o(intermediate_reg_2[607])); 
fsm fsm_inst_2_293(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1213]),.i2(intermediate_reg_1[1212]),.o(intermediate_reg_2[606])); 
mux_module mux_module_inst_2_294(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1211]),.i2(intermediate_reg_1[1210]),.o(intermediate_reg_2[605]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_295(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1209]),.i2(intermediate_reg_1[1208]),.o(intermediate_reg_2[604])); 
mux_module mux_module_inst_2_296(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1207]),.i2(intermediate_reg_1[1206]),.o(intermediate_reg_2[603]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_297(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1205]),.i2(intermediate_reg_1[1204]),.o(intermediate_reg_2[602])); 
mux_module mux_module_inst_2_298(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1203]),.i2(intermediate_reg_1[1202]),.o(intermediate_reg_2[601]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_299(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1201]),.i2(intermediate_reg_1[1200]),.o(intermediate_reg_2[600])); 
mux_module mux_module_inst_2_300(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1199]),.i2(intermediate_reg_1[1198]),.o(intermediate_reg_2[599]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_301(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1197]),.i2(intermediate_reg_1[1196]),.o(intermediate_reg_2[598]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_302(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1195]),.i2(intermediate_reg_1[1194]),.o(intermediate_reg_2[597]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_303(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1193]),.i2(intermediate_reg_1[1192]),.o(intermediate_reg_2[596]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_304(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1191]),.i2(intermediate_reg_1[1190]),.o(intermediate_reg_2[595])); 
fsm fsm_inst_2_305(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1189]),.i2(intermediate_reg_1[1188]),.o(intermediate_reg_2[594])); 
fsm fsm_inst_2_306(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1187]),.i2(intermediate_reg_1[1186]),.o(intermediate_reg_2[593])); 
mux_module mux_module_inst_2_307(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1185]),.i2(intermediate_reg_1[1184]),.o(intermediate_reg_2[592]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_308(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1183]),.i2(intermediate_reg_1[1182]),.o(intermediate_reg_2[591])); 
mux_module mux_module_inst_2_309(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1181]),.i2(intermediate_reg_1[1180]),.o(intermediate_reg_2[590]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_310(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1179]),.i2(intermediate_reg_1[1178]),.o(intermediate_reg_2[589])); 
fsm fsm_inst_2_311(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1177]),.i2(intermediate_reg_1[1176]),.o(intermediate_reg_2[588])); 
mux_module mux_module_inst_2_312(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1175]),.i2(intermediate_reg_1[1174]),.o(intermediate_reg_2[587]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_313(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1173]),.i2(intermediate_reg_1[1172]),.o(intermediate_reg_2[586])); 
fsm fsm_inst_2_314(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1171]),.i2(intermediate_reg_1[1170]),.o(intermediate_reg_2[585])); 
fsm fsm_inst_2_315(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1169]),.i2(intermediate_reg_1[1168]),.o(intermediate_reg_2[584])); 
mux_module mux_module_inst_2_316(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1167]),.i2(intermediate_reg_1[1166]),.o(intermediate_reg_2[583]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_317(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1165]),.i2(intermediate_reg_1[1164]),.o(intermediate_reg_2[582])); 
fsm fsm_inst_2_318(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1163]),.i2(intermediate_reg_1[1162]),.o(intermediate_reg_2[581])); 
mux_module mux_module_inst_2_319(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1161]),.i2(intermediate_reg_1[1160]),.o(intermediate_reg_2[580]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_320(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1159]),.i2(intermediate_reg_1[1158]),.o(intermediate_reg_2[579]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_321(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1157]),.i2(intermediate_reg_1[1156]),.o(intermediate_reg_2[578]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_322(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1155]),.i2(intermediate_reg_1[1154]),.o(intermediate_reg_2[577]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_323(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1153]),.i2(intermediate_reg_1[1152]),.o(intermediate_reg_2[576]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_324(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1151]),.i2(intermediate_reg_1[1150]),.o(intermediate_reg_2[575])); 
mux_module mux_module_inst_2_325(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1149]),.i2(intermediate_reg_1[1148]),.o(intermediate_reg_2[574]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_326(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1147]),.i2(intermediate_reg_1[1146]),.o(intermediate_reg_2[573])); 
fsm fsm_inst_2_327(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1145]),.i2(intermediate_reg_1[1144]),.o(intermediate_reg_2[572])); 
fsm fsm_inst_2_328(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1143]),.i2(intermediate_reg_1[1142]),.o(intermediate_reg_2[571])); 
mux_module mux_module_inst_2_329(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1141]),.i2(intermediate_reg_1[1140]),.o(intermediate_reg_2[570]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_330(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1139]),.i2(intermediate_reg_1[1138]),.o(intermediate_reg_2[569]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_331(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1137]),.i2(intermediate_reg_1[1136]),.o(intermediate_reg_2[568])); 
fsm fsm_inst_2_332(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1135]),.i2(intermediate_reg_1[1134]),.o(intermediate_reg_2[567])); 
mux_module mux_module_inst_2_333(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1133]),.i2(intermediate_reg_1[1132]),.o(intermediate_reg_2[566]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_334(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1131]),.i2(intermediate_reg_1[1130]),.o(intermediate_reg_2[565])); 
mux_module mux_module_inst_2_335(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1129]),.i2(intermediate_reg_1[1128]),.o(intermediate_reg_2[564]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_336(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1127]),.i2(intermediate_reg_1[1126]),.o(intermediate_reg_2[563])); 
fsm fsm_inst_2_337(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1125]),.i2(intermediate_reg_1[1124]),.o(intermediate_reg_2[562])); 
fsm fsm_inst_2_338(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1123]),.i2(intermediate_reg_1[1122]),.o(intermediate_reg_2[561])); 
fsm fsm_inst_2_339(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1121]),.i2(intermediate_reg_1[1120]),.o(intermediate_reg_2[560])); 
fsm fsm_inst_2_340(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1119]),.i2(intermediate_reg_1[1118]),.o(intermediate_reg_2[559])); 
mux_module mux_module_inst_2_341(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1117]),.i2(intermediate_reg_1[1116]),.o(intermediate_reg_2[558]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_342(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1115]),.i2(intermediate_reg_1[1114]),.o(intermediate_reg_2[557])); 
fsm fsm_inst_2_343(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1113]),.i2(intermediate_reg_1[1112]),.o(intermediate_reg_2[556])); 
fsm fsm_inst_2_344(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1111]),.i2(intermediate_reg_1[1110]),.o(intermediate_reg_2[555])); 
fsm fsm_inst_2_345(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1109]),.i2(intermediate_reg_1[1108]),.o(intermediate_reg_2[554])); 
mux_module mux_module_inst_2_346(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1107]),.i2(intermediate_reg_1[1106]),.o(intermediate_reg_2[553]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_347(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1105]),.i2(intermediate_reg_1[1104]),.o(intermediate_reg_2[552])); 
mux_module mux_module_inst_2_348(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1103]),.i2(intermediate_reg_1[1102]),.o(intermediate_reg_2[551]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_349(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1101]),.i2(intermediate_reg_1[1100]),.o(intermediate_reg_2[550])); 
mux_module mux_module_inst_2_350(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1099]),.i2(intermediate_reg_1[1098]),.o(intermediate_reg_2[549]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_351(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1097]),.i2(intermediate_reg_1[1096]),.o(intermediate_reg_2[548]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_352(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1095]),.i2(intermediate_reg_1[1094]),.o(intermediate_reg_2[547]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_353(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1093]),.i2(intermediate_reg_1[1092]),.o(intermediate_reg_2[546]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_354(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1091]),.i2(intermediate_reg_1[1090]),.o(intermediate_reg_2[545]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_355(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1089]),.i2(intermediate_reg_1[1088]),.o(intermediate_reg_2[544])); 
mux_module mux_module_inst_2_356(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1087]),.i2(intermediate_reg_1[1086]),.o(intermediate_reg_2[543]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_357(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1085]),.i2(intermediate_reg_1[1084]),.o(intermediate_reg_2[542]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_358(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1083]),.i2(intermediate_reg_1[1082]),.o(intermediate_reg_2[541]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_359(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1081]),.i2(intermediate_reg_1[1080]),.o(intermediate_reg_2[540]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_360(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1079]),.i2(intermediate_reg_1[1078]),.o(intermediate_reg_2[539])); 
mux_module mux_module_inst_2_361(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1077]),.i2(intermediate_reg_1[1076]),.o(intermediate_reg_2[538]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_362(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1075]),.i2(intermediate_reg_1[1074]),.o(intermediate_reg_2[537])); 
fsm fsm_inst_2_363(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1073]),.i2(intermediate_reg_1[1072]),.o(intermediate_reg_2[536])); 
fsm fsm_inst_2_364(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1071]),.i2(intermediate_reg_1[1070]),.o(intermediate_reg_2[535])); 
fsm fsm_inst_2_365(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1069]),.i2(intermediate_reg_1[1068]),.o(intermediate_reg_2[534])); 
mux_module mux_module_inst_2_366(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1067]),.i2(intermediate_reg_1[1066]),.o(intermediate_reg_2[533]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_367(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1065]),.i2(intermediate_reg_1[1064]),.o(intermediate_reg_2[532]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_368(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1063]),.i2(intermediate_reg_1[1062]),.o(intermediate_reg_2[531]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_369(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1061]),.i2(intermediate_reg_1[1060]),.o(intermediate_reg_2[530]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_370(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1059]),.i2(intermediate_reg_1[1058]),.o(intermediate_reg_2[529])); 
mux_module mux_module_inst_2_371(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1057]),.i2(intermediate_reg_1[1056]),.o(intermediate_reg_2[528]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_372(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1055]),.i2(intermediate_reg_1[1054]),.o(intermediate_reg_2[527])); 
fsm fsm_inst_2_373(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1053]),.i2(intermediate_reg_1[1052]),.o(intermediate_reg_2[526])); 
mux_module mux_module_inst_2_374(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1051]),.i2(intermediate_reg_1[1050]),.o(intermediate_reg_2[525]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_375(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1049]),.i2(intermediate_reg_1[1048]),.o(intermediate_reg_2[524])); 
mux_module mux_module_inst_2_376(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1047]),.i2(intermediate_reg_1[1046]),.o(intermediate_reg_2[523]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_377(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1045]),.i2(intermediate_reg_1[1044]),.o(intermediate_reg_2[522]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_378(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1043]),.i2(intermediate_reg_1[1042]),.o(intermediate_reg_2[521]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_379(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1041]),.i2(intermediate_reg_1[1040]),.o(intermediate_reg_2[520]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_380(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1039]),.i2(intermediate_reg_1[1038]),.o(intermediate_reg_2[519]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_381(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1037]),.i2(intermediate_reg_1[1036]),.o(intermediate_reg_2[518])); 
mux_module mux_module_inst_2_382(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1035]),.i2(intermediate_reg_1[1034]),.o(intermediate_reg_2[517]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_383(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1033]),.i2(intermediate_reg_1[1032]),.o(intermediate_reg_2[516]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_384(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1031]),.i2(intermediate_reg_1[1030]),.o(intermediate_reg_2[515]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_385(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1029]),.i2(intermediate_reg_1[1028]),.o(intermediate_reg_2[514])); 
mux_module mux_module_inst_2_386(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1027]),.i2(intermediate_reg_1[1026]),.o(intermediate_reg_2[513]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_387(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1025]),.i2(intermediate_reg_1[1024]),.o(intermediate_reg_2[512]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_388(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1023]),.i2(intermediate_reg_1[1022]),.o(intermediate_reg_2[511]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_389(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1021]),.i2(intermediate_reg_1[1020]),.o(intermediate_reg_2[510])); 
fsm fsm_inst_2_390(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1019]),.i2(intermediate_reg_1[1018]),.o(intermediate_reg_2[509])); 
mux_module mux_module_inst_2_391(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1017]),.i2(intermediate_reg_1[1016]),.o(intermediate_reg_2[508]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_392(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1015]),.i2(intermediate_reg_1[1014]),.o(intermediate_reg_2[507])); 
fsm fsm_inst_2_393(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1013]),.i2(intermediate_reg_1[1012]),.o(intermediate_reg_2[506])); 
mux_module mux_module_inst_2_394(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1011]),.i2(intermediate_reg_1[1010]),.o(intermediate_reg_2[505]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_395(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1009]),.i2(intermediate_reg_1[1008]),.o(intermediate_reg_2[504])); 
fsm fsm_inst_2_396(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1007]),.i2(intermediate_reg_1[1006]),.o(intermediate_reg_2[503])); 
fsm fsm_inst_2_397(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1005]),.i2(intermediate_reg_1[1004]),.o(intermediate_reg_2[502])); 
fsm fsm_inst_2_398(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1003]),.i2(intermediate_reg_1[1002]),.o(intermediate_reg_2[501])); 
mux_module mux_module_inst_2_399(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1001]),.i2(intermediate_reg_1[1000]),.o(intermediate_reg_2[500]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_400(.clk(clk),.reset(reset),.i1(intermediate_reg_1[999]),.i2(intermediate_reg_1[998]),.o(intermediate_reg_2[499]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_401(.clk(clk),.reset(reset),.i1(intermediate_reg_1[997]),.i2(intermediate_reg_1[996]),.o(intermediate_reg_2[498]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_402(.clk(clk),.reset(reset),.i1(intermediate_reg_1[995]),.i2(intermediate_reg_1[994]),.o(intermediate_reg_2[497])); 
fsm fsm_inst_2_403(.clk(clk),.reset(reset),.i1(intermediate_reg_1[993]),.i2(intermediate_reg_1[992]),.o(intermediate_reg_2[496])); 
mux_module mux_module_inst_2_404(.clk(clk),.reset(reset),.i1(intermediate_reg_1[991]),.i2(intermediate_reg_1[990]),.o(intermediate_reg_2[495]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_405(.clk(clk),.reset(reset),.i1(intermediate_reg_1[989]),.i2(intermediate_reg_1[988]),.o(intermediate_reg_2[494])); 
fsm fsm_inst_2_406(.clk(clk),.reset(reset),.i1(intermediate_reg_1[987]),.i2(intermediate_reg_1[986]),.o(intermediate_reg_2[493])); 
mux_module mux_module_inst_2_407(.clk(clk),.reset(reset),.i1(intermediate_reg_1[985]),.i2(intermediate_reg_1[984]),.o(intermediate_reg_2[492]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_408(.clk(clk),.reset(reset),.i1(intermediate_reg_1[983]),.i2(intermediate_reg_1[982]),.o(intermediate_reg_2[491])); 
fsm fsm_inst_2_409(.clk(clk),.reset(reset),.i1(intermediate_reg_1[981]),.i2(intermediate_reg_1[980]),.o(intermediate_reg_2[490])); 
mux_module mux_module_inst_2_410(.clk(clk),.reset(reset),.i1(intermediate_reg_1[979]),.i2(intermediate_reg_1[978]),.o(intermediate_reg_2[489]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_411(.clk(clk),.reset(reset),.i1(intermediate_reg_1[977]),.i2(intermediate_reg_1[976]),.o(intermediate_reg_2[488])); 
fsm fsm_inst_2_412(.clk(clk),.reset(reset),.i1(intermediate_reg_1[975]),.i2(intermediate_reg_1[974]),.o(intermediate_reg_2[487])); 
mux_module mux_module_inst_2_413(.clk(clk),.reset(reset),.i1(intermediate_reg_1[973]),.i2(intermediate_reg_1[972]),.o(intermediate_reg_2[486]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_414(.clk(clk),.reset(reset),.i1(intermediate_reg_1[971]),.i2(intermediate_reg_1[970]),.o(intermediate_reg_2[485]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_415(.clk(clk),.reset(reset),.i1(intermediate_reg_1[969]),.i2(intermediate_reg_1[968]),.o(intermediate_reg_2[484]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_416(.clk(clk),.reset(reset),.i1(intermediate_reg_1[967]),.i2(intermediate_reg_1[966]),.o(intermediate_reg_2[483])); 
mux_module mux_module_inst_2_417(.clk(clk),.reset(reset),.i1(intermediate_reg_1[965]),.i2(intermediate_reg_1[964]),.o(intermediate_reg_2[482]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_418(.clk(clk),.reset(reset),.i1(intermediate_reg_1[963]),.i2(intermediate_reg_1[962]),.o(intermediate_reg_2[481]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_419(.clk(clk),.reset(reset),.i1(intermediate_reg_1[961]),.i2(intermediate_reg_1[960]),.o(intermediate_reg_2[480])); 
fsm fsm_inst_2_420(.clk(clk),.reset(reset),.i1(intermediate_reg_1[959]),.i2(intermediate_reg_1[958]),.o(intermediate_reg_2[479])); 
fsm fsm_inst_2_421(.clk(clk),.reset(reset),.i1(intermediate_reg_1[957]),.i2(intermediate_reg_1[956]),.o(intermediate_reg_2[478])); 
fsm fsm_inst_2_422(.clk(clk),.reset(reset),.i1(intermediate_reg_1[955]),.i2(intermediate_reg_1[954]),.o(intermediate_reg_2[477])); 
mux_module mux_module_inst_2_423(.clk(clk),.reset(reset),.i1(intermediate_reg_1[953]),.i2(intermediate_reg_1[952]),.o(intermediate_reg_2[476]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_424(.clk(clk),.reset(reset),.i1(intermediate_reg_1[951]),.i2(intermediate_reg_1[950]),.o(intermediate_reg_2[475])); 
mux_module mux_module_inst_2_425(.clk(clk),.reset(reset),.i1(intermediate_reg_1[949]),.i2(intermediate_reg_1[948]),.o(intermediate_reg_2[474]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_426(.clk(clk),.reset(reset),.i1(intermediate_reg_1[947]),.i2(intermediate_reg_1[946]),.o(intermediate_reg_2[473]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_427(.clk(clk),.reset(reset),.i1(intermediate_reg_1[945]),.i2(intermediate_reg_1[944]),.o(intermediate_reg_2[472])); 
fsm fsm_inst_2_428(.clk(clk),.reset(reset),.i1(intermediate_reg_1[943]),.i2(intermediate_reg_1[942]),.o(intermediate_reg_2[471])); 
fsm fsm_inst_2_429(.clk(clk),.reset(reset),.i1(intermediate_reg_1[941]),.i2(intermediate_reg_1[940]),.o(intermediate_reg_2[470])); 
mux_module mux_module_inst_2_430(.clk(clk),.reset(reset),.i1(intermediate_reg_1[939]),.i2(intermediate_reg_1[938]),.o(intermediate_reg_2[469]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_431(.clk(clk),.reset(reset),.i1(intermediate_reg_1[937]),.i2(intermediate_reg_1[936]),.o(intermediate_reg_2[468]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_432(.clk(clk),.reset(reset),.i1(intermediate_reg_1[935]),.i2(intermediate_reg_1[934]),.o(intermediate_reg_2[467]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_433(.clk(clk),.reset(reset),.i1(intermediate_reg_1[933]),.i2(intermediate_reg_1[932]),.o(intermediate_reg_2[466]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_434(.clk(clk),.reset(reset),.i1(intermediate_reg_1[931]),.i2(intermediate_reg_1[930]),.o(intermediate_reg_2[465]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_435(.clk(clk),.reset(reset),.i1(intermediate_reg_1[929]),.i2(intermediate_reg_1[928]),.o(intermediate_reg_2[464])); 
fsm fsm_inst_2_436(.clk(clk),.reset(reset),.i1(intermediate_reg_1[927]),.i2(intermediate_reg_1[926]),.o(intermediate_reg_2[463])); 
fsm fsm_inst_2_437(.clk(clk),.reset(reset),.i1(intermediate_reg_1[925]),.i2(intermediate_reg_1[924]),.o(intermediate_reg_2[462])); 
fsm fsm_inst_2_438(.clk(clk),.reset(reset),.i1(intermediate_reg_1[923]),.i2(intermediate_reg_1[922]),.o(intermediate_reg_2[461])); 
mux_module mux_module_inst_2_439(.clk(clk),.reset(reset),.i1(intermediate_reg_1[921]),.i2(intermediate_reg_1[920]),.o(intermediate_reg_2[460]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_440(.clk(clk),.reset(reset),.i1(intermediate_reg_1[919]),.i2(intermediate_reg_1[918]),.o(intermediate_reg_2[459])); 
mux_module mux_module_inst_2_441(.clk(clk),.reset(reset),.i1(intermediate_reg_1[917]),.i2(intermediate_reg_1[916]),.o(intermediate_reg_2[458]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_442(.clk(clk),.reset(reset),.i1(intermediate_reg_1[915]),.i2(intermediate_reg_1[914]),.o(intermediate_reg_2[457])); 
fsm fsm_inst_2_443(.clk(clk),.reset(reset),.i1(intermediate_reg_1[913]),.i2(intermediate_reg_1[912]),.o(intermediate_reg_2[456])); 
mux_module mux_module_inst_2_444(.clk(clk),.reset(reset),.i1(intermediate_reg_1[911]),.i2(intermediate_reg_1[910]),.o(intermediate_reg_2[455]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_445(.clk(clk),.reset(reset),.i1(intermediate_reg_1[909]),.i2(intermediate_reg_1[908]),.o(intermediate_reg_2[454])); 
mux_module mux_module_inst_2_446(.clk(clk),.reset(reset),.i1(intermediate_reg_1[907]),.i2(intermediate_reg_1[906]),.o(intermediate_reg_2[453]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_447(.clk(clk),.reset(reset),.i1(intermediate_reg_1[905]),.i2(intermediate_reg_1[904]),.o(intermediate_reg_2[452]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_448(.clk(clk),.reset(reset),.i1(intermediate_reg_1[903]),.i2(intermediate_reg_1[902]),.o(intermediate_reg_2[451]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_449(.clk(clk),.reset(reset),.i1(intermediate_reg_1[901]),.i2(intermediate_reg_1[900]),.o(intermediate_reg_2[450])); 
fsm fsm_inst_2_450(.clk(clk),.reset(reset),.i1(intermediate_reg_1[899]),.i2(intermediate_reg_1[898]),.o(intermediate_reg_2[449])); 
mux_module mux_module_inst_2_451(.clk(clk),.reset(reset),.i1(intermediate_reg_1[897]),.i2(intermediate_reg_1[896]),.o(intermediate_reg_2[448]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_452(.clk(clk),.reset(reset),.i1(intermediate_reg_1[895]),.i2(intermediate_reg_1[894]),.o(intermediate_reg_2[447])); 
mux_module mux_module_inst_2_453(.clk(clk),.reset(reset),.i1(intermediate_reg_1[893]),.i2(intermediate_reg_1[892]),.o(intermediate_reg_2[446]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_454(.clk(clk),.reset(reset),.i1(intermediate_reg_1[891]),.i2(intermediate_reg_1[890]),.o(intermediate_reg_2[445])); 
mux_module mux_module_inst_2_455(.clk(clk),.reset(reset),.i1(intermediate_reg_1[889]),.i2(intermediate_reg_1[888]),.o(intermediate_reg_2[444]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_456(.clk(clk),.reset(reset),.i1(intermediate_reg_1[887]),.i2(intermediate_reg_1[886]),.o(intermediate_reg_2[443]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_457(.clk(clk),.reset(reset),.i1(intermediate_reg_1[885]),.i2(intermediate_reg_1[884]),.o(intermediate_reg_2[442])); 
fsm fsm_inst_2_458(.clk(clk),.reset(reset),.i1(intermediate_reg_1[883]),.i2(intermediate_reg_1[882]),.o(intermediate_reg_2[441])); 
mux_module mux_module_inst_2_459(.clk(clk),.reset(reset),.i1(intermediate_reg_1[881]),.i2(intermediate_reg_1[880]),.o(intermediate_reg_2[440]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_460(.clk(clk),.reset(reset),.i1(intermediate_reg_1[879]),.i2(intermediate_reg_1[878]),.o(intermediate_reg_2[439])); 
mux_module mux_module_inst_2_461(.clk(clk),.reset(reset),.i1(intermediate_reg_1[877]),.i2(intermediate_reg_1[876]),.o(intermediate_reg_2[438]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_462(.clk(clk),.reset(reset),.i1(intermediate_reg_1[875]),.i2(intermediate_reg_1[874]),.o(intermediate_reg_2[437])); 
mux_module mux_module_inst_2_463(.clk(clk),.reset(reset),.i1(intermediate_reg_1[873]),.i2(intermediate_reg_1[872]),.o(intermediate_reg_2[436]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_464(.clk(clk),.reset(reset),.i1(intermediate_reg_1[871]),.i2(intermediate_reg_1[870]),.o(intermediate_reg_2[435]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_465(.clk(clk),.reset(reset),.i1(intermediate_reg_1[869]),.i2(intermediate_reg_1[868]),.o(intermediate_reg_2[434])); 
fsm fsm_inst_2_466(.clk(clk),.reset(reset),.i1(intermediate_reg_1[867]),.i2(intermediate_reg_1[866]),.o(intermediate_reg_2[433])); 
fsm fsm_inst_2_467(.clk(clk),.reset(reset),.i1(intermediate_reg_1[865]),.i2(intermediate_reg_1[864]),.o(intermediate_reg_2[432])); 
fsm fsm_inst_2_468(.clk(clk),.reset(reset),.i1(intermediate_reg_1[863]),.i2(intermediate_reg_1[862]),.o(intermediate_reg_2[431])); 
mux_module mux_module_inst_2_469(.clk(clk),.reset(reset),.i1(intermediate_reg_1[861]),.i2(intermediate_reg_1[860]),.o(intermediate_reg_2[430]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_470(.clk(clk),.reset(reset),.i1(intermediate_reg_1[859]),.i2(intermediate_reg_1[858]),.o(intermediate_reg_2[429])); 
mux_module mux_module_inst_2_471(.clk(clk),.reset(reset),.i1(intermediate_reg_1[857]),.i2(intermediate_reg_1[856]),.o(intermediate_reg_2[428]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_472(.clk(clk),.reset(reset),.i1(intermediate_reg_1[855]),.i2(intermediate_reg_1[854]),.o(intermediate_reg_2[427])); 
fsm fsm_inst_2_473(.clk(clk),.reset(reset),.i1(intermediate_reg_1[853]),.i2(intermediate_reg_1[852]),.o(intermediate_reg_2[426])); 
mux_module mux_module_inst_2_474(.clk(clk),.reset(reset),.i1(intermediate_reg_1[851]),.i2(intermediate_reg_1[850]),.o(intermediate_reg_2[425]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_475(.clk(clk),.reset(reset),.i1(intermediate_reg_1[849]),.i2(intermediate_reg_1[848]),.o(intermediate_reg_2[424]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_476(.clk(clk),.reset(reset),.i1(intermediate_reg_1[847]),.i2(intermediate_reg_1[846]),.o(intermediate_reg_2[423])); 
mux_module mux_module_inst_2_477(.clk(clk),.reset(reset),.i1(intermediate_reg_1[845]),.i2(intermediate_reg_1[844]),.o(intermediate_reg_2[422]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_478(.clk(clk),.reset(reset),.i1(intermediate_reg_1[843]),.i2(intermediate_reg_1[842]),.o(intermediate_reg_2[421]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_479(.clk(clk),.reset(reset),.i1(intermediate_reg_1[841]),.i2(intermediate_reg_1[840]),.o(intermediate_reg_2[420]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_480(.clk(clk),.reset(reset),.i1(intermediate_reg_1[839]),.i2(intermediate_reg_1[838]),.o(intermediate_reg_2[419])); 
fsm fsm_inst_2_481(.clk(clk),.reset(reset),.i1(intermediate_reg_1[837]),.i2(intermediate_reg_1[836]),.o(intermediate_reg_2[418])); 
fsm fsm_inst_2_482(.clk(clk),.reset(reset),.i1(intermediate_reg_1[835]),.i2(intermediate_reg_1[834]),.o(intermediate_reg_2[417])); 
fsm fsm_inst_2_483(.clk(clk),.reset(reset),.i1(intermediate_reg_1[833]),.i2(intermediate_reg_1[832]),.o(intermediate_reg_2[416])); 
mux_module mux_module_inst_2_484(.clk(clk),.reset(reset),.i1(intermediate_reg_1[831]),.i2(intermediate_reg_1[830]),.o(intermediate_reg_2[415]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_485(.clk(clk),.reset(reset),.i1(intermediate_reg_1[829]),.i2(intermediate_reg_1[828]),.o(intermediate_reg_2[414])); 
fsm fsm_inst_2_486(.clk(clk),.reset(reset),.i1(intermediate_reg_1[827]),.i2(intermediate_reg_1[826]),.o(intermediate_reg_2[413])); 
fsm fsm_inst_2_487(.clk(clk),.reset(reset),.i1(intermediate_reg_1[825]),.i2(intermediate_reg_1[824]),.o(intermediate_reg_2[412])); 
fsm fsm_inst_2_488(.clk(clk),.reset(reset),.i1(intermediate_reg_1[823]),.i2(intermediate_reg_1[822]),.o(intermediate_reg_2[411])); 
fsm fsm_inst_2_489(.clk(clk),.reset(reset),.i1(intermediate_reg_1[821]),.i2(intermediate_reg_1[820]),.o(intermediate_reg_2[410])); 
mux_module mux_module_inst_2_490(.clk(clk),.reset(reset),.i1(intermediate_reg_1[819]),.i2(intermediate_reg_1[818]),.o(intermediate_reg_2[409]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_491(.clk(clk),.reset(reset),.i1(intermediate_reg_1[817]),.i2(intermediate_reg_1[816]),.o(intermediate_reg_2[408])); 
fsm fsm_inst_2_492(.clk(clk),.reset(reset),.i1(intermediate_reg_1[815]),.i2(intermediate_reg_1[814]),.o(intermediate_reg_2[407])); 
fsm fsm_inst_2_493(.clk(clk),.reset(reset),.i1(intermediate_reg_1[813]),.i2(intermediate_reg_1[812]),.o(intermediate_reg_2[406])); 
mux_module mux_module_inst_2_494(.clk(clk),.reset(reset),.i1(intermediate_reg_1[811]),.i2(intermediate_reg_1[810]),.o(intermediate_reg_2[405]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_495(.clk(clk),.reset(reset),.i1(intermediate_reg_1[809]),.i2(intermediate_reg_1[808]),.o(intermediate_reg_2[404]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_496(.clk(clk),.reset(reset),.i1(intermediate_reg_1[807]),.i2(intermediate_reg_1[806]),.o(intermediate_reg_2[403])); 
mux_module mux_module_inst_2_497(.clk(clk),.reset(reset),.i1(intermediate_reg_1[805]),.i2(intermediate_reg_1[804]),.o(intermediate_reg_2[402]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_498(.clk(clk),.reset(reset),.i1(intermediate_reg_1[803]),.i2(intermediate_reg_1[802]),.o(intermediate_reg_2[401])); 
fsm fsm_inst_2_499(.clk(clk),.reset(reset),.i1(intermediate_reg_1[801]),.i2(intermediate_reg_1[800]),.o(intermediate_reg_2[400])); 
fsm fsm_inst_2_500(.clk(clk),.reset(reset),.i1(intermediate_reg_1[799]),.i2(intermediate_reg_1[798]),.o(intermediate_reg_2[399])); 
mux_module mux_module_inst_2_501(.clk(clk),.reset(reset),.i1(intermediate_reg_1[797]),.i2(intermediate_reg_1[796]),.o(intermediate_reg_2[398]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_502(.clk(clk),.reset(reset),.i1(intermediate_reg_1[795]),.i2(intermediate_reg_1[794]),.o(intermediate_reg_2[397])); 
mux_module mux_module_inst_2_503(.clk(clk),.reset(reset),.i1(intermediate_reg_1[793]),.i2(intermediate_reg_1[792]),.o(intermediate_reg_2[396]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_504(.clk(clk),.reset(reset),.i1(intermediate_reg_1[791]),.i2(intermediate_reg_1[790]),.o(intermediate_reg_2[395]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_505(.clk(clk),.reset(reset),.i1(intermediate_reg_1[789]),.i2(intermediate_reg_1[788]),.o(intermediate_reg_2[394]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_506(.clk(clk),.reset(reset),.i1(intermediate_reg_1[787]),.i2(intermediate_reg_1[786]),.o(intermediate_reg_2[393]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_507(.clk(clk),.reset(reset),.i1(intermediate_reg_1[785]),.i2(intermediate_reg_1[784]),.o(intermediate_reg_2[392]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_508(.clk(clk),.reset(reset),.i1(intermediate_reg_1[783]),.i2(intermediate_reg_1[782]),.o(intermediate_reg_2[391]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_509(.clk(clk),.reset(reset),.i1(intermediate_reg_1[781]),.i2(intermediate_reg_1[780]),.o(intermediate_reg_2[390]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_510(.clk(clk),.reset(reset),.i1(intermediate_reg_1[779]),.i2(intermediate_reg_1[778]),.o(intermediate_reg_2[389]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_511(.clk(clk),.reset(reset),.i1(intermediate_reg_1[777]),.i2(intermediate_reg_1[776]),.o(intermediate_reg_2[388])); 
mux_module mux_module_inst_2_512(.clk(clk),.reset(reset),.i1(intermediate_reg_1[775]),.i2(intermediate_reg_1[774]),.o(intermediate_reg_2[387]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_513(.clk(clk),.reset(reset),.i1(intermediate_reg_1[773]),.i2(intermediate_reg_1[772]),.o(intermediate_reg_2[386])); 
mux_module mux_module_inst_2_514(.clk(clk),.reset(reset),.i1(intermediate_reg_1[771]),.i2(intermediate_reg_1[770]),.o(intermediate_reg_2[385]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_515(.clk(clk),.reset(reset),.i1(intermediate_reg_1[769]),.i2(intermediate_reg_1[768]),.o(intermediate_reg_2[384]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_516(.clk(clk),.reset(reset),.i1(intermediate_reg_1[767]),.i2(intermediate_reg_1[766]),.o(intermediate_reg_2[383]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_517(.clk(clk),.reset(reset),.i1(intermediate_reg_1[765]),.i2(intermediate_reg_1[764]),.o(intermediate_reg_2[382]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_518(.clk(clk),.reset(reset),.i1(intermediate_reg_1[763]),.i2(intermediate_reg_1[762]),.o(intermediate_reg_2[381])); 
fsm fsm_inst_2_519(.clk(clk),.reset(reset),.i1(intermediate_reg_1[761]),.i2(intermediate_reg_1[760]),.o(intermediate_reg_2[380])); 
fsm fsm_inst_2_520(.clk(clk),.reset(reset),.i1(intermediate_reg_1[759]),.i2(intermediate_reg_1[758]),.o(intermediate_reg_2[379])); 
mux_module mux_module_inst_2_521(.clk(clk),.reset(reset),.i1(intermediate_reg_1[757]),.i2(intermediate_reg_1[756]),.o(intermediate_reg_2[378]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_522(.clk(clk),.reset(reset),.i1(intermediate_reg_1[755]),.i2(intermediate_reg_1[754]),.o(intermediate_reg_2[377])); 
fsm fsm_inst_2_523(.clk(clk),.reset(reset),.i1(intermediate_reg_1[753]),.i2(intermediate_reg_1[752]),.o(intermediate_reg_2[376])); 
fsm fsm_inst_2_524(.clk(clk),.reset(reset),.i1(intermediate_reg_1[751]),.i2(intermediate_reg_1[750]),.o(intermediate_reg_2[375])); 
mux_module mux_module_inst_2_525(.clk(clk),.reset(reset),.i1(intermediate_reg_1[749]),.i2(intermediate_reg_1[748]),.o(intermediate_reg_2[374]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_526(.clk(clk),.reset(reset),.i1(intermediate_reg_1[747]),.i2(intermediate_reg_1[746]),.o(intermediate_reg_2[373]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_527(.clk(clk),.reset(reset),.i1(intermediate_reg_1[745]),.i2(intermediate_reg_1[744]),.o(intermediate_reg_2[372])); 
mux_module mux_module_inst_2_528(.clk(clk),.reset(reset),.i1(intermediate_reg_1[743]),.i2(intermediate_reg_1[742]),.o(intermediate_reg_2[371]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_529(.clk(clk),.reset(reset),.i1(intermediate_reg_1[741]),.i2(intermediate_reg_1[740]),.o(intermediate_reg_2[370]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_530(.clk(clk),.reset(reset),.i1(intermediate_reg_1[739]),.i2(intermediate_reg_1[738]),.o(intermediate_reg_2[369]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_531(.clk(clk),.reset(reset),.i1(intermediate_reg_1[737]),.i2(intermediate_reg_1[736]),.o(intermediate_reg_2[368]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_532(.clk(clk),.reset(reset),.i1(intermediate_reg_1[735]),.i2(intermediate_reg_1[734]),.o(intermediate_reg_2[367]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_533(.clk(clk),.reset(reset),.i1(intermediate_reg_1[733]),.i2(intermediate_reg_1[732]),.o(intermediate_reg_2[366]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_534(.clk(clk),.reset(reset),.i1(intermediate_reg_1[731]),.i2(intermediate_reg_1[730]),.o(intermediate_reg_2[365]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_535(.clk(clk),.reset(reset),.i1(intermediate_reg_1[729]),.i2(intermediate_reg_1[728]),.o(intermediate_reg_2[364]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_536(.clk(clk),.reset(reset),.i1(intermediate_reg_1[727]),.i2(intermediate_reg_1[726]),.o(intermediate_reg_2[363])); 
fsm fsm_inst_2_537(.clk(clk),.reset(reset),.i1(intermediate_reg_1[725]),.i2(intermediate_reg_1[724]),.o(intermediate_reg_2[362])); 
fsm fsm_inst_2_538(.clk(clk),.reset(reset),.i1(intermediate_reg_1[723]),.i2(intermediate_reg_1[722]),.o(intermediate_reg_2[361])); 
mux_module mux_module_inst_2_539(.clk(clk),.reset(reset),.i1(intermediate_reg_1[721]),.i2(intermediate_reg_1[720]),.o(intermediate_reg_2[360]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_540(.clk(clk),.reset(reset),.i1(intermediate_reg_1[719]),.i2(intermediate_reg_1[718]),.o(intermediate_reg_2[359]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_541(.clk(clk),.reset(reset),.i1(intermediate_reg_1[717]),.i2(intermediate_reg_1[716]),.o(intermediate_reg_2[358])); 
fsm fsm_inst_2_542(.clk(clk),.reset(reset),.i1(intermediate_reg_1[715]),.i2(intermediate_reg_1[714]),.o(intermediate_reg_2[357])); 
fsm fsm_inst_2_543(.clk(clk),.reset(reset),.i1(intermediate_reg_1[713]),.i2(intermediate_reg_1[712]),.o(intermediate_reg_2[356])); 
fsm fsm_inst_2_544(.clk(clk),.reset(reset),.i1(intermediate_reg_1[711]),.i2(intermediate_reg_1[710]),.o(intermediate_reg_2[355])); 
mux_module mux_module_inst_2_545(.clk(clk),.reset(reset),.i1(intermediate_reg_1[709]),.i2(intermediate_reg_1[708]),.o(intermediate_reg_2[354]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_546(.clk(clk),.reset(reset),.i1(intermediate_reg_1[707]),.i2(intermediate_reg_1[706]),.o(intermediate_reg_2[353])); 
mux_module mux_module_inst_2_547(.clk(clk),.reset(reset),.i1(intermediate_reg_1[705]),.i2(intermediate_reg_1[704]),.o(intermediate_reg_2[352]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_548(.clk(clk),.reset(reset),.i1(intermediate_reg_1[703]),.i2(intermediate_reg_1[702]),.o(intermediate_reg_2[351]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_549(.clk(clk),.reset(reset),.i1(intermediate_reg_1[701]),.i2(intermediate_reg_1[700]),.o(intermediate_reg_2[350]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_550(.clk(clk),.reset(reset),.i1(intermediate_reg_1[699]),.i2(intermediate_reg_1[698]),.o(intermediate_reg_2[349])); 
mux_module mux_module_inst_2_551(.clk(clk),.reset(reset),.i1(intermediate_reg_1[697]),.i2(intermediate_reg_1[696]),.o(intermediate_reg_2[348]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_552(.clk(clk),.reset(reset),.i1(intermediate_reg_1[695]),.i2(intermediate_reg_1[694]),.o(intermediate_reg_2[347])); 
fsm fsm_inst_2_553(.clk(clk),.reset(reset),.i1(intermediate_reg_1[693]),.i2(intermediate_reg_1[692]),.o(intermediate_reg_2[346])); 
mux_module mux_module_inst_2_554(.clk(clk),.reset(reset),.i1(intermediate_reg_1[691]),.i2(intermediate_reg_1[690]),.o(intermediate_reg_2[345]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_555(.clk(clk),.reset(reset),.i1(intermediate_reg_1[689]),.i2(intermediate_reg_1[688]),.o(intermediate_reg_2[344])); 
mux_module mux_module_inst_2_556(.clk(clk),.reset(reset),.i1(intermediate_reg_1[687]),.i2(intermediate_reg_1[686]),.o(intermediate_reg_2[343]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_557(.clk(clk),.reset(reset),.i1(intermediate_reg_1[685]),.i2(intermediate_reg_1[684]),.o(intermediate_reg_2[342]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_558(.clk(clk),.reset(reset),.i1(intermediate_reg_1[683]),.i2(intermediate_reg_1[682]),.o(intermediate_reg_2[341])); 
fsm fsm_inst_2_559(.clk(clk),.reset(reset),.i1(intermediate_reg_1[681]),.i2(intermediate_reg_1[680]),.o(intermediate_reg_2[340])); 
mux_module mux_module_inst_2_560(.clk(clk),.reset(reset),.i1(intermediate_reg_1[679]),.i2(intermediate_reg_1[678]),.o(intermediate_reg_2[339]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_561(.clk(clk),.reset(reset),.i1(intermediate_reg_1[677]),.i2(intermediate_reg_1[676]),.o(intermediate_reg_2[338]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_562(.clk(clk),.reset(reset),.i1(intermediate_reg_1[675]),.i2(intermediate_reg_1[674]),.o(intermediate_reg_2[337])); 
mux_module mux_module_inst_2_563(.clk(clk),.reset(reset),.i1(intermediate_reg_1[673]),.i2(intermediate_reg_1[672]),.o(intermediate_reg_2[336]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_564(.clk(clk),.reset(reset),.i1(intermediate_reg_1[671]),.i2(intermediate_reg_1[670]),.o(intermediate_reg_2[335])); 
mux_module mux_module_inst_2_565(.clk(clk),.reset(reset),.i1(intermediate_reg_1[669]),.i2(intermediate_reg_1[668]),.o(intermediate_reg_2[334]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_566(.clk(clk),.reset(reset),.i1(intermediate_reg_1[667]),.i2(intermediate_reg_1[666]),.o(intermediate_reg_2[333]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_567(.clk(clk),.reset(reset),.i1(intermediate_reg_1[665]),.i2(intermediate_reg_1[664]),.o(intermediate_reg_2[332])); 
mux_module mux_module_inst_2_568(.clk(clk),.reset(reset),.i1(intermediate_reg_1[663]),.i2(intermediate_reg_1[662]),.o(intermediate_reg_2[331]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_569(.clk(clk),.reset(reset),.i1(intermediate_reg_1[661]),.i2(intermediate_reg_1[660]),.o(intermediate_reg_2[330]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_570(.clk(clk),.reset(reset),.i1(intermediate_reg_1[659]),.i2(intermediate_reg_1[658]),.o(intermediate_reg_2[329])); 
fsm fsm_inst_2_571(.clk(clk),.reset(reset),.i1(intermediate_reg_1[657]),.i2(intermediate_reg_1[656]),.o(intermediate_reg_2[328])); 
mux_module mux_module_inst_2_572(.clk(clk),.reset(reset),.i1(intermediate_reg_1[655]),.i2(intermediate_reg_1[654]),.o(intermediate_reg_2[327]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_573(.clk(clk),.reset(reset),.i1(intermediate_reg_1[653]),.i2(intermediate_reg_1[652]),.o(intermediate_reg_2[326]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_574(.clk(clk),.reset(reset),.i1(intermediate_reg_1[651]),.i2(intermediate_reg_1[650]),.o(intermediate_reg_2[325])); 
mux_module mux_module_inst_2_575(.clk(clk),.reset(reset),.i1(intermediate_reg_1[649]),.i2(intermediate_reg_1[648]),.o(intermediate_reg_2[324]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_576(.clk(clk),.reset(reset),.i1(intermediate_reg_1[647]),.i2(intermediate_reg_1[646]),.o(intermediate_reg_2[323]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_577(.clk(clk),.reset(reset),.i1(intermediate_reg_1[645]),.i2(intermediate_reg_1[644]),.o(intermediate_reg_2[322])); 
mux_module mux_module_inst_2_578(.clk(clk),.reset(reset),.i1(intermediate_reg_1[643]),.i2(intermediate_reg_1[642]),.o(intermediate_reg_2[321]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_579(.clk(clk),.reset(reset),.i1(intermediate_reg_1[641]),.i2(intermediate_reg_1[640]),.o(intermediate_reg_2[320]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_580(.clk(clk),.reset(reset),.i1(intermediate_reg_1[639]),.i2(intermediate_reg_1[638]),.o(intermediate_reg_2[319]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_581(.clk(clk),.reset(reset),.i1(intermediate_reg_1[637]),.i2(intermediate_reg_1[636]),.o(intermediate_reg_2[318])); 
fsm fsm_inst_2_582(.clk(clk),.reset(reset),.i1(intermediate_reg_1[635]),.i2(intermediate_reg_1[634]),.o(intermediate_reg_2[317])); 
fsm fsm_inst_2_583(.clk(clk),.reset(reset),.i1(intermediate_reg_1[633]),.i2(intermediate_reg_1[632]),.o(intermediate_reg_2[316])); 
fsm fsm_inst_2_584(.clk(clk),.reset(reset),.i1(intermediate_reg_1[631]),.i2(intermediate_reg_1[630]),.o(intermediate_reg_2[315])); 
mux_module mux_module_inst_2_585(.clk(clk),.reset(reset),.i1(intermediate_reg_1[629]),.i2(intermediate_reg_1[628]),.o(intermediate_reg_2[314]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_586(.clk(clk),.reset(reset),.i1(intermediate_reg_1[627]),.i2(intermediate_reg_1[626]),.o(intermediate_reg_2[313]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_587(.clk(clk),.reset(reset),.i1(intermediate_reg_1[625]),.i2(intermediate_reg_1[624]),.o(intermediate_reg_2[312])); 
fsm fsm_inst_2_588(.clk(clk),.reset(reset),.i1(intermediate_reg_1[623]),.i2(intermediate_reg_1[622]),.o(intermediate_reg_2[311])); 
mux_module mux_module_inst_2_589(.clk(clk),.reset(reset),.i1(intermediate_reg_1[621]),.i2(intermediate_reg_1[620]),.o(intermediate_reg_2[310]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_590(.clk(clk),.reset(reset),.i1(intermediate_reg_1[619]),.i2(intermediate_reg_1[618]),.o(intermediate_reg_2[309])); 
fsm fsm_inst_2_591(.clk(clk),.reset(reset),.i1(intermediate_reg_1[617]),.i2(intermediate_reg_1[616]),.o(intermediate_reg_2[308])); 
mux_module mux_module_inst_2_592(.clk(clk),.reset(reset),.i1(intermediate_reg_1[615]),.i2(intermediate_reg_1[614]),.o(intermediate_reg_2[307]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_593(.clk(clk),.reset(reset),.i1(intermediate_reg_1[613]),.i2(intermediate_reg_1[612]),.o(intermediate_reg_2[306]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_594(.clk(clk),.reset(reset),.i1(intermediate_reg_1[611]),.i2(intermediate_reg_1[610]),.o(intermediate_reg_2[305])); 
fsm fsm_inst_2_595(.clk(clk),.reset(reset),.i1(intermediate_reg_1[609]),.i2(intermediate_reg_1[608]),.o(intermediate_reg_2[304])); 
fsm fsm_inst_2_596(.clk(clk),.reset(reset),.i1(intermediate_reg_1[607]),.i2(intermediate_reg_1[606]),.o(intermediate_reg_2[303])); 
mux_module mux_module_inst_2_597(.clk(clk),.reset(reset),.i1(intermediate_reg_1[605]),.i2(intermediate_reg_1[604]),.o(intermediate_reg_2[302]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_598(.clk(clk),.reset(reset),.i1(intermediate_reg_1[603]),.i2(intermediate_reg_1[602]),.o(intermediate_reg_2[301])); 
fsm fsm_inst_2_599(.clk(clk),.reset(reset),.i1(intermediate_reg_1[601]),.i2(intermediate_reg_1[600]),.o(intermediate_reg_2[300])); 
fsm fsm_inst_2_600(.clk(clk),.reset(reset),.i1(intermediate_reg_1[599]),.i2(intermediate_reg_1[598]),.o(intermediate_reg_2[299])); 
fsm fsm_inst_2_601(.clk(clk),.reset(reset),.i1(intermediate_reg_1[597]),.i2(intermediate_reg_1[596]),.o(intermediate_reg_2[298])); 
mux_module mux_module_inst_2_602(.clk(clk),.reset(reset),.i1(intermediate_reg_1[595]),.i2(intermediate_reg_1[594]),.o(intermediate_reg_2[297]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_603(.clk(clk),.reset(reset),.i1(intermediate_reg_1[593]),.i2(intermediate_reg_1[592]),.o(intermediate_reg_2[296])); 
fsm fsm_inst_2_604(.clk(clk),.reset(reset),.i1(intermediate_reg_1[591]),.i2(intermediate_reg_1[590]),.o(intermediate_reg_2[295])); 
mux_module mux_module_inst_2_605(.clk(clk),.reset(reset),.i1(intermediate_reg_1[589]),.i2(intermediate_reg_1[588]),.o(intermediate_reg_2[294]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_606(.clk(clk),.reset(reset),.i1(intermediate_reg_1[587]),.i2(intermediate_reg_1[586]),.o(intermediate_reg_2[293])); 
fsm fsm_inst_2_607(.clk(clk),.reset(reset),.i1(intermediate_reg_1[585]),.i2(intermediate_reg_1[584]),.o(intermediate_reg_2[292])); 
fsm fsm_inst_2_608(.clk(clk),.reset(reset),.i1(intermediate_reg_1[583]),.i2(intermediate_reg_1[582]),.o(intermediate_reg_2[291])); 
mux_module mux_module_inst_2_609(.clk(clk),.reset(reset),.i1(intermediate_reg_1[581]),.i2(intermediate_reg_1[580]),.o(intermediate_reg_2[290]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_610(.clk(clk),.reset(reset),.i1(intermediate_reg_1[579]),.i2(intermediate_reg_1[578]),.o(intermediate_reg_2[289]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_611(.clk(clk),.reset(reset),.i1(intermediate_reg_1[577]),.i2(intermediate_reg_1[576]),.o(intermediate_reg_2[288]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_612(.clk(clk),.reset(reset),.i1(intermediate_reg_1[575]),.i2(intermediate_reg_1[574]),.o(intermediate_reg_2[287])); 
mux_module mux_module_inst_2_613(.clk(clk),.reset(reset),.i1(intermediate_reg_1[573]),.i2(intermediate_reg_1[572]),.o(intermediate_reg_2[286]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_614(.clk(clk),.reset(reset),.i1(intermediate_reg_1[571]),.i2(intermediate_reg_1[570]),.o(intermediate_reg_2[285]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_615(.clk(clk),.reset(reset),.i1(intermediate_reg_1[569]),.i2(intermediate_reg_1[568]),.o(intermediate_reg_2[284])); 
mux_module mux_module_inst_2_616(.clk(clk),.reset(reset),.i1(intermediate_reg_1[567]),.i2(intermediate_reg_1[566]),.o(intermediate_reg_2[283]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_617(.clk(clk),.reset(reset),.i1(intermediate_reg_1[565]),.i2(intermediate_reg_1[564]),.o(intermediate_reg_2[282]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_618(.clk(clk),.reset(reset),.i1(intermediate_reg_1[563]),.i2(intermediate_reg_1[562]),.o(intermediate_reg_2[281]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_619(.clk(clk),.reset(reset),.i1(intermediate_reg_1[561]),.i2(intermediate_reg_1[560]),.o(intermediate_reg_2[280])); 
mux_module mux_module_inst_2_620(.clk(clk),.reset(reset),.i1(intermediate_reg_1[559]),.i2(intermediate_reg_1[558]),.o(intermediate_reg_2[279]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_621(.clk(clk),.reset(reset),.i1(intermediate_reg_1[557]),.i2(intermediate_reg_1[556]),.o(intermediate_reg_2[278]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_622(.clk(clk),.reset(reset),.i1(intermediate_reg_1[555]),.i2(intermediate_reg_1[554]),.o(intermediate_reg_2[277]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_623(.clk(clk),.reset(reset),.i1(intermediate_reg_1[553]),.i2(intermediate_reg_1[552]),.o(intermediate_reg_2[276])); 
fsm fsm_inst_2_624(.clk(clk),.reset(reset),.i1(intermediate_reg_1[551]),.i2(intermediate_reg_1[550]),.o(intermediate_reg_2[275])); 
mux_module mux_module_inst_2_625(.clk(clk),.reset(reset),.i1(intermediate_reg_1[549]),.i2(intermediate_reg_1[548]),.o(intermediate_reg_2[274]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_626(.clk(clk),.reset(reset),.i1(intermediate_reg_1[547]),.i2(intermediate_reg_1[546]),.o(intermediate_reg_2[273])); 
fsm fsm_inst_2_627(.clk(clk),.reset(reset),.i1(intermediate_reg_1[545]),.i2(intermediate_reg_1[544]),.o(intermediate_reg_2[272])); 
fsm fsm_inst_2_628(.clk(clk),.reset(reset),.i1(intermediate_reg_1[543]),.i2(intermediate_reg_1[542]),.o(intermediate_reg_2[271])); 
mux_module mux_module_inst_2_629(.clk(clk),.reset(reset),.i1(intermediate_reg_1[541]),.i2(intermediate_reg_1[540]),.o(intermediate_reg_2[270]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_630(.clk(clk),.reset(reset),.i1(intermediate_reg_1[539]),.i2(intermediate_reg_1[538]),.o(intermediate_reg_2[269]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_631(.clk(clk),.reset(reset),.i1(intermediate_reg_1[537]),.i2(intermediate_reg_1[536]),.o(intermediate_reg_2[268])); 
mux_module mux_module_inst_2_632(.clk(clk),.reset(reset),.i1(intermediate_reg_1[535]),.i2(intermediate_reg_1[534]),.o(intermediate_reg_2[267]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_633(.clk(clk),.reset(reset),.i1(intermediate_reg_1[533]),.i2(intermediate_reg_1[532]),.o(intermediate_reg_2[266])); 
mux_module mux_module_inst_2_634(.clk(clk),.reset(reset),.i1(intermediate_reg_1[531]),.i2(intermediate_reg_1[530]),.o(intermediate_reg_2[265]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_635(.clk(clk),.reset(reset),.i1(intermediate_reg_1[529]),.i2(intermediate_reg_1[528]),.o(intermediate_reg_2[264]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_636(.clk(clk),.reset(reset),.i1(intermediate_reg_1[527]),.i2(intermediate_reg_1[526]),.o(intermediate_reg_2[263]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_637(.clk(clk),.reset(reset),.i1(intermediate_reg_1[525]),.i2(intermediate_reg_1[524]),.o(intermediate_reg_2[262])); 
mux_module mux_module_inst_2_638(.clk(clk),.reset(reset),.i1(intermediate_reg_1[523]),.i2(intermediate_reg_1[522]),.o(intermediate_reg_2[261]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_639(.clk(clk),.reset(reset),.i1(intermediate_reg_1[521]),.i2(intermediate_reg_1[520]),.o(intermediate_reg_2[260])); 
fsm fsm_inst_2_640(.clk(clk),.reset(reset),.i1(intermediate_reg_1[519]),.i2(intermediate_reg_1[518]),.o(intermediate_reg_2[259])); 
fsm fsm_inst_2_641(.clk(clk),.reset(reset),.i1(intermediate_reg_1[517]),.i2(intermediate_reg_1[516]),.o(intermediate_reg_2[258])); 
fsm fsm_inst_2_642(.clk(clk),.reset(reset),.i1(intermediate_reg_1[515]),.i2(intermediate_reg_1[514]),.o(intermediate_reg_2[257])); 
fsm fsm_inst_2_643(.clk(clk),.reset(reset),.i1(intermediate_reg_1[513]),.i2(intermediate_reg_1[512]),.o(intermediate_reg_2[256])); 
fsm fsm_inst_2_644(.clk(clk),.reset(reset),.i1(intermediate_reg_1[511]),.i2(intermediate_reg_1[510]),.o(intermediate_reg_2[255])); 
mux_module mux_module_inst_2_645(.clk(clk),.reset(reset),.i1(intermediate_reg_1[509]),.i2(intermediate_reg_1[508]),.o(intermediate_reg_2[254]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_646(.clk(clk),.reset(reset),.i1(intermediate_reg_1[507]),.i2(intermediate_reg_1[506]),.o(intermediate_reg_2[253])); 
mux_module mux_module_inst_2_647(.clk(clk),.reset(reset),.i1(intermediate_reg_1[505]),.i2(intermediate_reg_1[504]),.o(intermediate_reg_2[252]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_648(.clk(clk),.reset(reset),.i1(intermediate_reg_1[503]),.i2(intermediate_reg_1[502]),.o(intermediate_reg_2[251])); 
fsm fsm_inst_2_649(.clk(clk),.reset(reset),.i1(intermediate_reg_1[501]),.i2(intermediate_reg_1[500]),.o(intermediate_reg_2[250])); 
fsm fsm_inst_2_650(.clk(clk),.reset(reset),.i1(intermediate_reg_1[499]),.i2(intermediate_reg_1[498]),.o(intermediate_reg_2[249])); 
mux_module mux_module_inst_2_651(.clk(clk),.reset(reset),.i1(intermediate_reg_1[497]),.i2(intermediate_reg_1[496]),.o(intermediate_reg_2[248]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_652(.clk(clk),.reset(reset),.i1(intermediate_reg_1[495]),.i2(intermediate_reg_1[494]),.o(intermediate_reg_2[247]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_653(.clk(clk),.reset(reset),.i1(intermediate_reg_1[493]),.i2(intermediate_reg_1[492]),.o(intermediate_reg_2[246]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_654(.clk(clk),.reset(reset),.i1(intermediate_reg_1[491]),.i2(intermediate_reg_1[490]),.o(intermediate_reg_2[245])); 
mux_module mux_module_inst_2_655(.clk(clk),.reset(reset),.i1(intermediate_reg_1[489]),.i2(intermediate_reg_1[488]),.o(intermediate_reg_2[244]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_656(.clk(clk),.reset(reset),.i1(intermediate_reg_1[487]),.i2(intermediate_reg_1[486]),.o(intermediate_reg_2[243]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_657(.clk(clk),.reset(reset),.i1(intermediate_reg_1[485]),.i2(intermediate_reg_1[484]),.o(intermediate_reg_2[242])); 
mux_module mux_module_inst_2_658(.clk(clk),.reset(reset),.i1(intermediate_reg_1[483]),.i2(intermediate_reg_1[482]),.o(intermediate_reg_2[241]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_659(.clk(clk),.reset(reset),.i1(intermediate_reg_1[481]),.i2(intermediate_reg_1[480]),.o(intermediate_reg_2[240]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_660(.clk(clk),.reset(reset),.i1(intermediate_reg_1[479]),.i2(intermediate_reg_1[478]),.o(intermediate_reg_2[239])); 
fsm fsm_inst_2_661(.clk(clk),.reset(reset),.i1(intermediate_reg_1[477]),.i2(intermediate_reg_1[476]),.o(intermediate_reg_2[238])); 
fsm fsm_inst_2_662(.clk(clk),.reset(reset),.i1(intermediate_reg_1[475]),.i2(intermediate_reg_1[474]),.o(intermediate_reg_2[237])); 
fsm fsm_inst_2_663(.clk(clk),.reset(reset),.i1(intermediate_reg_1[473]),.i2(intermediate_reg_1[472]),.o(intermediate_reg_2[236])); 
fsm fsm_inst_2_664(.clk(clk),.reset(reset),.i1(intermediate_reg_1[471]),.i2(intermediate_reg_1[470]),.o(intermediate_reg_2[235])); 
mux_module mux_module_inst_2_665(.clk(clk),.reset(reset),.i1(intermediate_reg_1[469]),.i2(intermediate_reg_1[468]),.o(intermediate_reg_2[234]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_666(.clk(clk),.reset(reset),.i1(intermediate_reg_1[467]),.i2(intermediate_reg_1[466]),.o(intermediate_reg_2[233]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_667(.clk(clk),.reset(reset),.i1(intermediate_reg_1[465]),.i2(intermediate_reg_1[464]),.o(intermediate_reg_2[232]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_668(.clk(clk),.reset(reset),.i1(intermediate_reg_1[463]),.i2(intermediate_reg_1[462]),.o(intermediate_reg_2[231]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_669(.clk(clk),.reset(reset),.i1(intermediate_reg_1[461]),.i2(intermediate_reg_1[460]),.o(intermediate_reg_2[230]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_670(.clk(clk),.reset(reset),.i1(intermediate_reg_1[459]),.i2(intermediate_reg_1[458]),.o(intermediate_reg_2[229]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_671(.clk(clk),.reset(reset),.i1(intermediate_reg_1[457]),.i2(intermediate_reg_1[456]),.o(intermediate_reg_2[228])); 
mux_module mux_module_inst_2_672(.clk(clk),.reset(reset),.i1(intermediate_reg_1[455]),.i2(intermediate_reg_1[454]),.o(intermediate_reg_2[227]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_673(.clk(clk),.reset(reset),.i1(intermediate_reg_1[453]),.i2(intermediate_reg_1[452]),.o(intermediate_reg_2[226]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_674(.clk(clk),.reset(reset),.i1(intermediate_reg_1[451]),.i2(intermediate_reg_1[450]),.o(intermediate_reg_2[225])); 
fsm fsm_inst_2_675(.clk(clk),.reset(reset),.i1(intermediate_reg_1[449]),.i2(intermediate_reg_1[448]),.o(intermediate_reg_2[224])); 
mux_module mux_module_inst_2_676(.clk(clk),.reset(reset),.i1(intermediate_reg_1[447]),.i2(intermediate_reg_1[446]),.o(intermediate_reg_2[223]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_677(.clk(clk),.reset(reset),.i1(intermediate_reg_1[445]),.i2(intermediate_reg_1[444]),.o(intermediate_reg_2[222])); 
fsm fsm_inst_2_678(.clk(clk),.reset(reset),.i1(intermediate_reg_1[443]),.i2(intermediate_reg_1[442]),.o(intermediate_reg_2[221])); 
mux_module mux_module_inst_2_679(.clk(clk),.reset(reset),.i1(intermediate_reg_1[441]),.i2(intermediate_reg_1[440]),.o(intermediate_reg_2[220]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_680(.clk(clk),.reset(reset),.i1(intermediate_reg_1[439]),.i2(intermediate_reg_1[438]),.o(intermediate_reg_2[219])); 
mux_module mux_module_inst_2_681(.clk(clk),.reset(reset),.i1(intermediate_reg_1[437]),.i2(intermediate_reg_1[436]),.o(intermediate_reg_2[218]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_682(.clk(clk),.reset(reset),.i1(intermediate_reg_1[435]),.i2(intermediate_reg_1[434]),.o(intermediate_reg_2[217]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_683(.clk(clk),.reset(reset),.i1(intermediate_reg_1[433]),.i2(intermediate_reg_1[432]),.o(intermediate_reg_2[216]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_684(.clk(clk),.reset(reset),.i1(intermediate_reg_1[431]),.i2(intermediate_reg_1[430]),.o(intermediate_reg_2[215])); 
mux_module mux_module_inst_2_685(.clk(clk),.reset(reset),.i1(intermediate_reg_1[429]),.i2(intermediate_reg_1[428]),.o(intermediate_reg_2[214]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_686(.clk(clk),.reset(reset),.i1(intermediate_reg_1[427]),.i2(intermediate_reg_1[426]),.o(intermediate_reg_2[213])); 
fsm fsm_inst_2_687(.clk(clk),.reset(reset),.i1(intermediate_reg_1[425]),.i2(intermediate_reg_1[424]),.o(intermediate_reg_2[212])); 
fsm fsm_inst_2_688(.clk(clk),.reset(reset),.i1(intermediate_reg_1[423]),.i2(intermediate_reg_1[422]),.o(intermediate_reg_2[211])); 
mux_module mux_module_inst_2_689(.clk(clk),.reset(reset),.i1(intermediate_reg_1[421]),.i2(intermediate_reg_1[420]),.o(intermediate_reg_2[210]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_690(.clk(clk),.reset(reset),.i1(intermediate_reg_1[419]),.i2(intermediate_reg_1[418]),.o(intermediate_reg_2[209])); 
mux_module mux_module_inst_2_691(.clk(clk),.reset(reset),.i1(intermediate_reg_1[417]),.i2(intermediate_reg_1[416]),.o(intermediate_reg_2[208]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_692(.clk(clk),.reset(reset),.i1(intermediate_reg_1[415]),.i2(intermediate_reg_1[414]),.o(intermediate_reg_2[207])); 
fsm fsm_inst_2_693(.clk(clk),.reset(reset),.i1(intermediate_reg_1[413]),.i2(intermediate_reg_1[412]),.o(intermediate_reg_2[206])); 
fsm fsm_inst_2_694(.clk(clk),.reset(reset),.i1(intermediate_reg_1[411]),.i2(intermediate_reg_1[410]),.o(intermediate_reg_2[205])); 
fsm fsm_inst_2_695(.clk(clk),.reset(reset),.i1(intermediate_reg_1[409]),.i2(intermediate_reg_1[408]),.o(intermediate_reg_2[204])); 
fsm fsm_inst_2_696(.clk(clk),.reset(reset),.i1(intermediate_reg_1[407]),.i2(intermediate_reg_1[406]),.o(intermediate_reg_2[203])); 
fsm fsm_inst_2_697(.clk(clk),.reset(reset),.i1(intermediate_reg_1[405]),.i2(intermediate_reg_1[404]),.o(intermediate_reg_2[202])); 
fsm fsm_inst_2_698(.clk(clk),.reset(reset),.i1(intermediate_reg_1[403]),.i2(intermediate_reg_1[402]),.o(intermediate_reg_2[201])); 
mux_module mux_module_inst_2_699(.clk(clk),.reset(reset),.i1(intermediate_reg_1[401]),.i2(intermediate_reg_1[400]),.o(intermediate_reg_2[200]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_700(.clk(clk),.reset(reset),.i1(intermediate_reg_1[399]),.i2(intermediate_reg_1[398]),.o(intermediate_reg_2[199])); 
fsm fsm_inst_2_701(.clk(clk),.reset(reset),.i1(intermediate_reg_1[397]),.i2(intermediate_reg_1[396]),.o(intermediate_reg_2[198])); 
mux_module mux_module_inst_2_702(.clk(clk),.reset(reset),.i1(intermediate_reg_1[395]),.i2(intermediate_reg_1[394]),.o(intermediate_reg_2[197]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_703(.clk(clk),.reset(reset),.i1(intermediate_reg_1[393]),.i2(intermediate_reg_1[392]),.o(intermediate_reg_2[196])); 
mux_module mux_module_inst_2_704(.clk(clk),.reset(reset),.i1(intermediate_reg_1[391]),.i2(intermediate_reg_1[390]),.o(intermediate_reg_2[195]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_705(.clk(clk),.reset(reset),.i1(intermediate_reg_1[389]),.i2(intermediate_reg_1[388]),.o(intermediate_reg_2[194]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_706(.clk(clk),.reset(reset),.i1(intermediate_reg_1[387]),.i2(intermediate_reg_1[386]),.o(intermediate_reg_2[193]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_707(.clk(clk),.reset(reset),.i1(intermediate_reg_1[385]),.i2(intermediate_reg_1[384]),.o(intermediate_reg_2[192]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_708(.clk(clk),.reset(reset),.i1(intermediate_reg_1[383]),.i2(intermediate_reg_1[382]),.o(intermediate_reg_2[191]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_709(.clk(clk),.reset(reset),.i1(intermediate_reg_1[381]),.i2(intermediate_reg_1[380]),.o(intermediate_reg_2[190]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_710(.clk(clk),.reset(reset),.i1(intermediate_reg_1[379]),.i2(intermediate_reg_1[378]),.o(intermediate_reg_2[189])); 
fsm fsm_inst_2_711(.clk(clk),.reset(reset),.i1(intermediate_reg_1[377]),.i2(intermediate_reg_1[376]),.o(intermediate_reg_2[188])); 
mux_module mux_module_inst_2_712(.clk(clk),.reset(reset),.i1(intermediate_reg_1[375]),.i2(intermediate_reg_1[374]),.o(intermediate_reg_2[187]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_713(.clk(clk),.reset(reset),.i1(intermediate_reg_1[373]),.i2(intermediate_reg_1[372]),.o(intermediate_reg_2[186])); 
mux_module mux_module_inst_2_714(.clk(clk),.reset(reset),.i1(intermediate_reg_1[371]),.i2(intermediate_reg_1[370]),.o(intermediate_reg_2[185]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_715(.clk(clk),.reset(reset),.i1(intermediate_reg_1[369]),.i2(intermediate_reg_1[368]),.o(intermediate_reg_2[184]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_716(.clk(clk),.reset(reset),.i1(intermediate_reg_1[367]),.i2(intermediate_reg_1[366]),.o(intermediate_reg_2[183]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_717(.clk(clk),.reset(reset),.i1(intermediate_reg_1[365]),.i2(intermediate_reg_1[364]),.o(intermediate_reg_2[182]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_718(.clk(clk),.reset(reset),.i1(intermediate_reg_1[363]),.i2(intermediate_reg_1[362]),.o(intermediate_reg_2[181]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_719(.clk(clk),.reset(reset),.i1(intermediate_reg_1[361]),.i2(intermediate_reg_1[360]),.o(intermediate_reg_2[180]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_720(.clk(clk),.reset(reset),.i1(intermediate_reg_1[359]),.i2(intermediate_reg_1[358]),.o(intermediate_reg_2[179]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_721(.clk(clk),.reset(reset),.i1(intermediate_reg_1[357]),.i2(intermediate_reg_1[356]),.o(intermediate_reg_2[178]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_722(.clk(clk),.reset(reset),.i1(intermediate_reg_1[355]),.i2(intermediate_reg_1[354]),.o(intermediate_reg_2[177]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_723(.clk(clk),.reset(reset),.i1(intermediate_reg_1[353]),.i2(intermediate_reg_1[352]),.o(intermediate_reg_2[176])); 
mux_module mux_module_inst_2_724(.clk(clk),.reset(reset),.i1(intermediate_reg_1[351]),.i2(intermediate_reg_1[350]),.o(intermediate_reg_2[175]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_725(.clk(clk),.reset(reset),.i1(intermediate_reg_1[349]),.i2(intermediate_reg_1[348]),.o(intermediate_reg_2[174]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_726(.clk(clk),.reset(reset),.i1(intermediate_reg_1[347]),.i2(intermediate_reg_1[346]),.o(intermediate_reg_2[173])); 
mux_module mux_module_inst_2_727(.clk(clk),.reset(reset),.i1(intermediate_reg_1[345]),.i2(intermediate_reg_1[344]),.o(intermediate_reg_2[172]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_728(.clk(clk),.reset(reset),.i1(intermediate_reg_1[343]),.i2(intermediate_reg_1[342]),.o(intermediate_reg_2[171])); 
fsm fsm_inst_2_729(.clk(clk),.reset(reset),.i1(intermediate_reg_1[341]),.i2(intermediate_reg_1[340]),.o(intermediate_reg_2[170])); 
mux_module mux_module_inst_2_730(.clk(clk),.reset(reset),.i1(intermediate_reg_1[339]),.i2(intermediate_reg_1[338]),.o(intermediate_reg_2[169]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_731(.clk(clk),.reset(reset),.i1(intermediate_reg_1[337]),.i2(intermediate_reg_1[336]),.o(intermediate_reg_2[168]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_732(.clk(clk),.reset(reset),.i1(intermediate_reg_1[335]),.i2(intermediate_reg_1[334]),.o(intermediate_reg_2[167]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_733(.clk(clk),.reset(reset),.i1(intermediate_reg_1[333]),.i2(intermediate_reg_1[332]),.o(intermediate_reg_2[166]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_734(.clk(clk),.reset(reset),.i1(intermediate_reg_1[331]),.i2(intermediate_reg_1[330]),.o(intermediate_reg_2[165]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_735(.clk(clk),.reset(reset),.i1(intermediate_reg_1[329]),.i2(intermediate_reg_1[328]),.o(intermediate_reg_2[164]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_736(.clk(clk),.reset(reset),.i1(intermediate_reg_1[327]),.i2(intermediate_reg_1[326]),.o(intermediate_reg_2[163])); 
mux_module mux_module_inst_2_737(.clk(clk),.reset(reset),.i1(intermediate_reg_1[325]),.i2(intermediate_reg_1[324]),.o(intermediate_reg_2[162]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_738(.clk(clk),.reset(reset),.i1(intermediate_reg_1[323]),.i2(intermediate_reg_1[322]),.o(intermediate_reg_2[161])); 
mux_module mux_module_inst_2_739(.clk(clk),.reset(reset),.i1(intermediate_reg_1[321]),.i2(intermediate_reg_1[320]),.o(intermediate_reg_2[160]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_740(.clk(clk),.reset(reset),.i1(intermediate_reg_1[319]),.i2(intermediate_reg_1[318]),.o(intermediate_reg_2[159])); 
fsm fsm_inst_2_741(.clk(clk),.reset(reset),.i1(intermediate_reg_1[317]),.i2(intermediate_reg_1[316]),.o(intermediate_reg_2[158])); 
fsm fsm_inst_2_742(.clk(clk),.reset(reset),.i1(intermediate_reg_1[315]),.i2(intermediate_reg_1[314]),.o(intermediate_reg_2[157])); 
mux_module mux_module_inst_2_743(.clk(clk),.reset(reset),.i1(intermediate_reg_1[313]),.i2(intermediate_reg_1[312]),.o(intermediate_reg_2[156]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_744(.clk(clk),.reset(reset),.i1(intermediate_reg_1[311]),.i2(intermediate_reg_1[310]),.o(intermediate_reg_2[155])); 
fsm fsm_inst_2_745(.clk(clk),.reset(reset),.i1(intermediate_reg_1[309]),.i2(intermediate_reg_1[308]),.o(intermediate_reg_2[154])); 
mux_module mux_module_inst_2_746(.clk(clk),.reset(reset),.i1(intermediate_reg_1[307]),.i2(intermediate_reg_1[306]),.o(intermediate_reg_2[153]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_747(.clk(clk),.reset(reset),.i1(intermediate_reg_1[305]),.i2(intermediate_reg_1[304]),.o(intermediate_reg_2[152]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_748(.clk(clk),.reset(reset),.i1(intermediate_reg_1[303]),.i2(intermediate_reg_1[302]),.o(intermediate_reg_2[151]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_749(.clk(clk),.reset(reset),.i1(intermediate_reg_1[301]),.i2(intermediate_reg_1[300]),.o(intermediate_reg_2[150])); 
fsm fsm_inst_2_750(.clk(clk),.reset(reset),.i1(intermediate_reg_1[299]),.i2(intermediate_reg_1[298]),.o(intermediate_reg_2[149])); 
fsm fsm_inst_2_751(.clk(clk),.reset(reset),.i1(intermediate_reg_1[297]),.i2(intermediate_reg_1[296]),.o(intermediate_reg_2[148])); 
mux_module mux_module_inst_2_752(.clk(clk),.reset(reset),.i1(intermediate_reg_1[295]),.i2(intermediate_reg_1[294]),.o(intermediate_reg_2[147]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_753(.clk(clk),.reset(reset),.i1(intermediate_reg_1[293]),.i2(intermediate_reg_1[292]),.o(intermediate_reg_2[146]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_754(.clk(clk),.reset(reset),.i1(intermediate_reg_1[291]),.i2(intermediate_reg_1[290]),.o(intermediate_reg_2[145]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_755(.clk(clk),.reset(reset),.i1(intermediate_reg_1[289]),.i2(intermediate_reg_1[288]),.o(intermediate_reg_2[144]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_756(.clk(clk),.reset(reset),.i1(intermediate_reg_1[287]),.i2(intermediate_reg_1[286]),.o(intermediate_reg_2[143])); 
fsm fsm_inst_2_757(.clk(clk),.reset(reset),.i1(intermediate_reg_1[285]),.i2(intermediate_reg_1[284]),.o(intermediate_reg_2[142])); 
mux_module mux_module_inst_2_758(.clk(clk),.reset(reset),.i1(intermediate_reg_1[283]),.i2(intermediate_reg_1[282]),.o(intermediate_reg_2[141]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_759(.clk(clk),.reset(reset),.i1(intermediate_reg_1[281]),.i2(intermediate_reg_1[280]),.o(intermediate_reg_2[140]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_760(.clk(clk),.reset(reset),.i1(intermediate_reg_1[279]),.i2(intermediate_reg_1[278]),.o(intermediate_reg_2[139])); 
mux_module mux_module_inst_2_761(.clk(clk),.reset(reset),.i1(intermediate_reg_1[277]),.i2(intermediate_reg_1[276]),.o(intermediate_reg_2[138]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_762(.clk(clk),.reset(reset),.i1(intermediate_reg_1[275]),.i2(intermediate_reg_1[274]),.o(intermediate_reg_2[137])); 
fsm fsm_inst_2_763(.clk(clk),.reset(reset),.i1(intermediate_reg_1[273]),.i2(intermediate_reg_1[272]),.o(intermediate_reg_2[136])); 
fsm fsm_inst_2_764(.clk(clk),.reset(reset),.i1(intermediate_reg_1[271]),.i2(intermediate_reg_1[270]),.o(intermediate_reg_2[135])); 
fsm fsm_inst_2_765(.clk(clk),.reset(reset),.i1(intermediate_reg_1[269]),.i2(intermediate_reg_1[268]),.o(intermediate_reg_2[134])); 
fsm fsm_inst_2_766(.clk(clk),.reset(reset),.i1(intermediate_reg_1[267]),.i2(intermediate_reg_1[266]),.o(intermediate_reg_2[133])); 
mux_module mux_module_inst_2_767(.clk(clk),.reset(reset),.i1(intermediate_reg_1[265]),.i2(intermediate_reg_1[264]),.o(intermediate_reg_2[132]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_768(.clk(clk),.reset(reset),.i1(intermediate_reg_1[263]),.i2(intermediate_reg_1[262]),.o(intermediate_reg_2[131]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_769(.clk(clk),.reset(reset),.i1(intermediate_reg_1[261]),.i2(intermediate_reg_1[260]),.o(intermediate_reg_2[130])); 
mux_module mux_module_inst_2_770(.clk(clk),.reset(reset),.i1(intermediate_reg_1[259]),.i2(intermediate_reg_1[258]),.o(intermediate_reg_2[129]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_771(.clk(clk),.reset(reset),.i1(intermediate_reg_1[257]),.i2(intermediate_reg_1[256]),.o(intermediate_reg_2[128])); 
fsm fsm_inst_2_772(.clk(clk),.reset(reset),.i1(intermediate_reg_1[255]),.i2(intermediate_reg_1[254]),.o(intermediate_reg_2[127])); 
mux_module mux_module_inst_2_773(.clk(clk),.reset(reset),.i1(intermediate_reg_1[253]),.i2(intermediate_reg_1[252]),.o(intermediate_reg_2[126]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_774(.clk(clk),.reset(reset),.i1(intermediate_reg_1[251]),.i2(intermediate_reg_1[250]),.o(intermediate_reg_2[125])); 
mux_module mux_module_inst_2_775(.clk(clk),.reset(reset),.i1(intermediate_reg_1[249]),.i2(intermediate_reg_1[248]),.o(intermediate_reg_2[124]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_776(.clk(clk),.reset(reset),.i1(intermediate_reg_1[247]),.i2(intermediate_reg_1[246]),.o(intermediate_reg_2[123])); 
fsm fsm_inst_2_777(.clk(clk),.reset(reset),.i1(intermediate_reg_1[245]),.i2(intermediate_reg_1[244]),.o(intermediate_reg_2[122])); 
mux_module mux_module_inst_2_778(.clk(clk),.reset(reset),.i1(intermediate_reg_1[243]),.i2(intermediate_reg_1[242]),.o(intermediate_reg_2[121]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_779(.clk(clk),.reset(reset),.i1(intermediate_reg_1[241]),.i2(intermediate_reg_1[240]),.o(intermediate_reg_2[120])); 
mux_module mux_module_inst_2_780(.clk(clk),.reset(reset),.i1(intermediate_reg_1[239]),.i2(intermediate_reg_1[238]),.o(intermediate_reg_2[119]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_781(.clk(clk),.reset(reset),.i1(intermediate_reg_1[237]),.i2(intermediate_reg_1[236]),.o(intermediate_reg_2[118]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_782(.clk(clk),.reset(reset),.i1(intermediate_reg_1[235]),.i2(intermediate_reg_1[234]),.o(intermediate_reg_2[117])); 
mux_module mux_module_inst_2_783(.clk(clk),.reset(reset),.i1(intermediate_reg_1[233]),.i2(intermediate_reg_1[232]),.o(intermediate_reg_2[116]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_784(.clk(clk),.reset(reset),.i1(intermediate_reg_1[231]),.i2(intermediate_reg_1[230]),.o(intermediate_reg_2[115]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_785(.clk(clk),.reset(reset),.i1(intermediate_reg_1[229]),.i2(intermediate_reg_1[228]),.o(intermediate_reg_2[114])); 
mux_module mux_module_inst_2_786(.clk(clk),.reset(reset),.i1(intermediate_reg_1[227]),.i2(intermediate_reg_1[226]),.o(intermediate_reg_2[113]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_787(.clk(clk),.reset(reset),.i1(intermediate_reg_1[225]),.i2(intermediate_reg_1[224]),.o(intermediate_reg_2[112])); 
mux_module mux_module_inst_2_788(.clk(clk),.reset(reset),.i1(intermediate_reg_1[223]),.i2(intermediate_reg_1[222]),.o(intermediate_reg_2[111]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_789(.clk(clk),.reset(reset),.i1(intermediate_reg_1[221]),.i2(intermediate_reg_1[220]),.o(intermediate_reg_2[110]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_790(.clk(clk),.reset(reset),.i1(intermediate_reg_1[219]),.i2(intermediate_reg_1[218]),.o(intermediate_reg_2[109])); 
fsm fsm_inst_2_791(.clk(clk),.reset(reset),.i1(intermediate_reg_1[217]),.i2(intermediate_reg_1[216]),.o(intermediate_reg_2[108])); 
mux_module mux_module_inst_2_792(.clk(clk),.reset(reset),.i1(intermediate_reg_1[215]),.i2(intermediate_reg_1[214]),.o(intermediate_reg_2[107]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_793(.clk(clk),.reset(reset),.i1(intermediate_reg_1[213]),.i2(intermediate_reg_1[212]),.o(intermediate_reg_2[106])); 
mux_module mux_module_inst_2_794(.clk(clk),.reset(reset),.i1(intermediate_reg_1[211]),.i2(intermediate_reg_1[210]),.o(intermediate_reg_2[105]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_795(.clk(clk),.reset(reset),.i1(intermediate_reg_1[209]),.i2(intermediate_reg_1[208]),.o(intermediate_reg_2[104]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_796(.clk(clk),.reset(reset),.i1(intermediate_reg_1[207]),.i2(intermediate_reg_1[206]),.o(intermediate_reg_2[103]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_797(.clk(clk),.reset(reset),.i1(intermediate_reg_1[205]),.i2(intermediate_reg_1[204]),.o(intermediate_reg_2[102])); 
mux_module mux_module_inst_2_798(.clk(clk),.reset(reset),.i1(intermediate_reg_1[203]),.i2(intermediate_reg_1[202]),.o(intermediate_reg_2[101]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_799(.clk(clk),.reset(reset),.i1(intermediate_reg_1[201]),.i2(intermediate_reg_1[200]),.o(intermediate_reg_2[100]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_800(.clk(clk),.reset(reset),.i1(intermediate_reg_1[199]),.i2(intermediate_reg_1[198]),.o(intermediate_reg_2[99]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_801(.clk(clk),.reset(reset),.i1(intermediate_reg_1[197]),.i2(intermediate_reg_1[196]),.o(intermediate_reg_2[98]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_802(.clk(clk),.reset(reset),.i1(intermediate_reg_1[195]),.i2(intermediate_reg_1[194]),.o(intermediate_reg_2[97])); 
mux_module mux_module_inst_2_803(.clk(clk),.reset(reset),.i1(intermediate_reg_1[193]),.i2(intermediate_reg_1[192]),.o(intermediate_reg_2[96]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_804(.clk(clk),.reset(reset),.i1(intermediate_reg_1[191]),.i2(intermediate_reg_1[190]),.o(intermediate_reg_2[95]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_805(.clk(clk),.reset(reset),.i1(intermediate_reg_1[189]),.i2(intermediate_reg_1[188]),.o(intermediate_reg_2[94]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_806(.clk(clk),.reset(reset),.i1(intermediate_reg_1[187]),.i2(intermediate_reg_1[186]),.o(intermediate_reg_2[93])); 
fsm fsm_inst_2_807(.clk(clk),.reset(reset),.i1(intermediate_reg_1[185]),.i2(intermediate_reg_1[184]),.o(intermediate_reg_2[92])); 
mux_module mux_module_inst_2_808(.clk(clk),.reset(reset),.i1(intermediate_reg_1[183]),.i2(intermediate_reg_1[182]),.o(intermediate_reg_2[91]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_809(.clk(clk),.reset(reset),.i1(intermediate_reg_1[181]),.i2(intermediate_reg_1[180]),.o(intermediate_reg_2[90])); 
fsm fsm_inst_2_810(.clk(clk),.reset(reset),.i1(intermediate_reg_1[179]),.i2(intermediate_reg_1[178]),.o(intermediate_reg_2[89])); 
mux_module mux_module_inst_2_811(.clk(clk),.reset(reset),.i1(intermediate_reg_1[177]),.i2(intermediate_reg_1[176]),.o(intermediate_reg_2[88]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_812(.clk(clk),.reset(reset),.i1(intermediate_reg_1[175]),.i2(intermediate_reg_1[174]),.o(intermediate_reg_2[87])); 
fsm fsm_inst_2_813(.clk(clk),.reset(reset),.i1(intermediate_reg_1[173]),.i2(intermediate_reg_1[172]),.o(intermediate_reg_2[86])); 
mux_module mux_module_inst_2_814(.clk(clk),.reset(reset),.i1(intermediate_reg_1[171]),.i2(intermediate_reg_1[170]),.o(intermediate_reg_2[85]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_815(.clk(clk),.reset(reset),.i1(intermediate_reg_1[169]),.i2(intermediate_reg_1[168]),.o(intermediate_reg_2[84])); 
fsm fsm_inst_2_816(.clk(clk),.reset(reset),.i1(intermediate_reg_1[167]),.i2(intermediate_reg_1[166]),.o(intermediate_reg_2[83])); 
mux_module mux_module_inst_2_817(.clk(clk),.reset(reset),.i1(intermediate_reg_1[165]),.i2(intermediate_reg_1[164]),.o(intermediate_reg_2[82]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_818(.clk(clk),.reset(reset),.i1(intermediate_reg_1[163]),.i2(intermediate_reg_1[162]),.o(intermediate_reg_2[81]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_819(.clk(clk),.reset(reset),.i1(intermediate_reg_1[161]),.i2(intermediate_reg_1[160]),.o(intermediate_reg_2[80]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_820(.clk(clk),.reset(reset),.i1(intermediate_reg_1[159]),.i2(intermediate_reg_1[158]),.o(intermediate_reg_2[79]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_821(.clk(clk),.reset(reset),.i1(intermediate_reg_1[157]),.i2(intermediate_reg_1[156]),.o(intermediate_reg_2[78]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_822(.clk(clk),.reset(reset),.i1(intermediate_reg_1[155]),.i2(intermediate_reg_1[154]),.o(intermediate_reg_2[77]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_823(.clk(clk),.reset(reset),.i1(intermediate_reg_1[153]),.i2(intermediate_reg_1[152]),.o(intermediate_reg_2[76]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_824(.clk(clk),.reset(reset),.i1(intermediate_reg_1[151]),.i2(intermediate_reg_1[150]),.o(intermediate_reg_2[75])); 
mux_module mux_module_inst_2_825(.clk(clk),.reset(reset),.i1(intermediate_reg_1[149]),.i2(intermediate_reg_1[148]),.o(intermediate_reg_2[74]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_826(.clk(clk),.reset(reset),.i1(intermediate_reg_1[147]),.i2(intermediate_reg_1[146]),.o(intermediate_reg_2[73]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_827(.clk(clk),.reset(reset),.i1(intermediate_reg_1[145]),.i2(intermediate_reg_1[144]),.o(intermediate_reg_2[72]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_828(.clk(clk),.reset(reset),.i1(intermediate_reg_1[143]),.i2(intermediate_reg_1[142]),.o(intermediate_reg_2[71]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_829(.clk(clk),.reset(reset),.i1(intermediate_reg_1[141]),.i2(intermediate_reg_1[140]),.o(intermediate_reg_2[70]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_830(.clk(clk),.reset(reset),.i1(intermediate_reg_1[139]),.i2(intermediate_reg_1[138]),.o(intermediate_reg_2[69])); 
mux_module mux_module_inst_2_831(.clk(clk),.reset(reset),.i1(intermediate_reg_1[137]),.i2(intermediate_reg_1[136]),.o(intermediate_reg_2[68]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_832(.clk(clk),.reset(reset),.i1(intermediate_reg_1[135]),.i2(intermediate_reg_1[134]),.o(intermediate_reg_2[67])); 
mux_module mux_module_inst_2_833(.clk(clk),.reset(reset),.i1(intermediate_reg_1[133]),.i2(intermediate_reg_1[132]),.o(intermediate_reg_2[66]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_834(.clk(clk),.reset(reset),.i1(intermediate_reg_1[131]),.i2(intermediate_reg_1[130]),.o(intermediate_reg_2[65])); 
mux_module mux_module_inst_2_835(.clk(clk),.reset(reset),.i1(intermediate_reg_1[129]),.i2(intermediate_reg_1[128]),.o(intermediate_reg_2[64]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_836(.clk(clk),.reset(reset),.i1(intermediate_reg_1[127]),.i2(intermediate_reg_1[126]),.o(intermediate_reg_2[63]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_837(.clk(clk),.reset(reset),.i1(intermediate_reg_1[125]),.i2(intermediate_reg_1[124]),.o(intermediate_reg_2[62]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_838(.clk(clk),.reset(reset),.i1(intermediate_reg_1[123]),.i2(intermediate_reg_1[122]),.o(intermediate_reg_2[61])); 
fsm fsm_inst_2_839(.clk(clk),.reset(reset),.i1(intermediate_reg_1[121]),.i2(intermediate_reg_1[120]),.o(intermediate_reg_2[60])); 
mux_module mux_module_inst_2_840(.clk(clk),.reset(reset),.i1(intermediate_reg_1[119]),.i2(intermediate_reg_1[118]),.o(intermediate_reg_2[59]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_841(.clk(clk),.reset(reset),.i1(intermediate_reg_1[117]),.i2(intermediate_reg_1[116]),.o(intermediate_reg_2[58]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_842(.clk(clk),.reset(reset),.i1(intermediate_reg_1[115]),.i2(intermediate_reg_1[114]),.o(intermediate_reg_2[57])); 
mux_module mux_module_inst_2_843(.clk(clk),.reset(reset),.i1(intermediate_reg_1[113]),.i2(intermediate_reg_1[112]),.o(intermediate_reg_2[56]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_844(.clk(clk),.reset(reset),.i1(intermediate_reg_1[111]),.i2(intermediate_reg_1[110]),.o(intermediate_reg_2[55]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_845(.clk(clk),.reset(reset),.i1(intermediate_reg_1[109]),.i2(intermediate_reg_1[108]),.o(intermediate_reg_2[54])); 
fsm fsm_inst_2_846(.clk(clk),.reset(reset),.i1(intermediate_reg_1[107]),.i2(intermediate_reg_1[106]),.o(intermediate_reg_2[53])); 
fsm fsm_inst_2_847(.clk(clk),.reset(reset),.i1(intermediate_reg_1[105]),.i2(intermediate_reg_1[104]),.o(intermediate_reg_2[52])); 
mux_module mux_module_inst_2_848(.clk(clk),.reset(reset),.i1(intermediate_reg_1[103]),.i2(intermediate_reg_1[102]),.o(intermediate_reg_2[51]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_849(.clk(clk),.reset(reset),.i1(intermediate_reg_1[101]),.i2(intermediate_reg_1[100]),.o(intermediate_reg_2[50]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_850(.clk(clk),.reset(reset),.i1(intermediate_reg_1[99]),.i2(intermediate_reg_1[98]),.o(intermediate_reg_2[49])); 
mux_module mux_module_inst_2_851(.clk(clk),.reset(reset),.i1(intermediate_reg_1[97]),.i2(intermediate_reg_1[96]),.o(intermediate_reg_2[48]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_852(.clk(clk),.reset(reset),.i1(intermediate_reg_1[95]),.i2(intermediate_reg_1[94]),.o(intermediate_reg_2[47]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_853(.clk(clk),.reset(reset),.i1(intermediate_reg_1[93]),.i2(intermediate_reg_1[92]),.o(intermediate_reg_2[46])); 
fsm fsm_inst_2_854(.clk(clk),.reset(reset),.i1(intermediate_reg_1[91]),.i2(intermediate_reg_1[90]),.o(intermediate_reg_2[45])); 
mux_module mux_module_inst_2_855(.clk(clk),.reset(reset),.i1(intermediate_reg_1[89]),.i2(intermediate_reg_1[88]),.o(intermediate_reg_2[44]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_856(.clk(clk),.reset(reset),.i1(intermediate_reg_1[87]),.i2(intermediate_reg_1[86]),.o(intermediate_reg_2[43])); 
fsm fsm_inst_2_857(.clk(clk),.reset(reset),.i1(intermediate_reg_1[85]),.i2(intermediate_reg_1[84]),.o(intermediate_reg_2[42])); 
fsm fsm_inst_2_858(.clk(clk),.reset(reset),.i1(intermediate_reg_1[83]),.i2(intermediate_reg_1[82]),.o(intermediate_reg_2[41])); 
fsm fsm_inst_2_859(.clk(clk),.reset(reset),.i1(intermediate_reg_1[81]),.i2(intermediate_reg_1[80]),.o(intermediate_reg_2[40])); 
fsm fsm_inst_2_860(.clk(clk),.reset(reset),.i1(intermediate_reg_1[79]),.i2(intermediate_reg_1[78]),.o(intermediate_reg_2[39])); 
mux_module mux_module_inst_2_861(.clk(clk),.reset(reset),.i1(intermediate_reg_1[77]),.i2(intermediate_reg_1[76]),.o(intermediate_reg_2[38]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_862(.clk(clk),.reset(reset),.i1(intermediate_reg_1[75]),.i2(intermediate_reg_1[74]),.o(intermediate_reg_2[37])); 
mux_module mux_module_inst_2_863(.clk(clk),.reset(reset),.i1(intermediate_reg_1[73]),.i2(intermediate_reg_1[72]),.o(intermediate_reg_2[36]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_864(.clk(clk),.reset(reset),.i1(intermediate_reg_1[71]),.i2(intermediate_reg_1[70]),.o(intermediate_reg_2[35]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_865(.clk(clk),.reset(reset),.i1(intermediate_reg_1[69]),.i2(intermediate_reg_1[68]),.o(intermediate_reg_2[34])); 
mux_module mux_module_inst_2_866(.clk(clk),.reset(reset),.i1(intermediate_reg_1[67]),.i2(intermediate_reg_1[66]),.o(intermediate_reg_2[33]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_867(.clk(clk),.reset(reset),.i1(intermediate_reg_1[65]),.i2(intermediate_reg_1[64]),.o(intermediate_reg_2[32])); 
mux_module mux_module_inst_2_868(.clk(clk),.reset(reset),.i1(intermediate_reg_1[63]),.i2(intermediate_reg_1[62]),.o(intermediate_reg_2[31]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_869(.clk(clk),.reset(reset),.i1(intermediate_reg_1[61]),.i2(intermediate_reg_1[60]),.o(intermediate_reg_2[30])); 
fsm fsm_inst_2_870(.clk(clk),.reset(reset),.i1(intermediate_reg_1[59]),.i2(intermediate_reg_1[58]),.o(intermediate_reg_2[29])); 
fsm fsm_inst_2_871(.clk(clk),.reset(reset),.i1(intermediate_reg_1[57]),.i2(intermediate_reg_1[56]),.o(intermediate_reg_2[28])); 
mux_module mux_module_inst_2_872(.clk(clk),.reset(reset),.i1(intermediate_reg_1[55]),.i2(intermediate_reg_1[54]),.o(intermediate_reg_2[27]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_873(.clk(clk),.reset(reset),.i1(intermediate_reg_1[53]),.i2(intermediate_reg_1[52]),.o(intermediate_reg_2[26]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_874(.clk(clk),.reset(reset),.i1(intermediate_reg_1[51]),.i2(intermediate_reg_1[50]),.o(intermediate_reg_2[25])); 
mux_module mux_module_inst_2_875(.clk(clk),.reset(reset),.i1(intermediate_reg_1[49]),.i2(intermediate_reg_1[48]),.o(intermediate_reg_2[24]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_876(.clk(clk),.reset(reset),.i1(intermediate_reg_1[47]),.i2(intermediate_reg_1[46]),.o(intermediate_reg_2[23]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_877(.clk(clk),.reset(reset),.i1(intermediate_reg_1[45]),.i2(intermediate_reg_1[44]),.o(intermediate_reg_2[22]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_878(.clk(clk),.reset(reset),.i1(intermediate_reg_1[43]),.i2(intermediate_reg_1[42]),.o(intermediate_reg_2[21])); 
mux_module mux_module_inst_2_879(.clk(clk),.reset(reset),.i1(intermediate_reg_1[41]),.i2(intermediate_reg_1[40]),.o(intermediate_reg_2[20]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_880(.clk(clk),.reset(reset),.i1(intermediate_reg_1[39]),.i2(intermediate_reg_1[38]),.o(intermediate_reg_2[19])); 
fsm fsm_inst_2_881(.clk(clk),.reset(reset),.i1(intermediate_reg_1[37]),.i2(intermediate_reg_1[36]),.o(intermediate_reg_2[18])); 
mux_module mux_module_inst_2_882(.clk(clk),.reset(reset),.i1(intermediate_reg_1[35]),.i2(intermediate_reg_1[34]),.o(intermediate_reg_2[17]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_883(.clk(clk),.reset(reset),.i1(intermediate_reg_1[33]),.i2(intermediate_reg_1[32]),.o(intermediate_reg_2[16]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_884(.clk(clk),.reset(reset),.i1(intermediate_reg_1[31]),.i2(intermediate_reg_1[30]),.o(intermediate_reg_2[15]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_885(.clk(clk),.reset(reset),.i1(intermediate_reg_1[29]),.i2(intermediate_reg_1[28]),.o(intermediate_reg_2[14]),.sel(intermediate_reg_1[0])); 
mux_module mux_module_inst_2_886(.clk(clk),.reset(reset),.i1(intermediate_reg_1[27]),.i2(intermediate_reg_1[26]),.o(intermediate_reg_2[13]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_887(.clk(clk),.reset(reset),.i1(intermediate_reg_1[25]),.i2(intermediate_reg_1[24]),.o(intermediate_reg_2[12])); 
fsm fsm_inst_2_888(.clk(clk),.reset(reset),.i1(intermediate_reg_1[23]),.i2(intermediate_reg_1[22]),.o(intermediate_reg_2[11])); 
fsm fsm_inst_2_889(.clk(clk),.reset(reset),.i1(intermediate_reg_1[21]),.i2(intermediate_reg_1[20]),.o(intermediate_reg_2[10])); 
fsm fsm_inst_2_890(.clk(clk),.reset(reset),.i1(intermediate_reg_1[19]),.i2(intermediate_reg_1[18]),.o(intermediate_reg_2[9])); 
mux_module mux_module_inst_2_891(.clk(clk),.reset(reset),.i1(intermediate_reg_1[17]),.i2(intermediate_reg_1[16]),.o(intermediate_reg_2[8]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_892(.clk(clk),.reset(reset),.i1(intermediate_reg_1[15]),.i2(intermediate_reg_1[14]),.o(intermediate_reg_2[7])); 
mux_module mux_module_inst_2_893(.clk(clk),.reset(reset),.i1(intermediate_reg_1[13]),.i2(intermediate_reg_1[12]),.o(intermediate_reg_2[6]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_894(.clk(clk),.reset(reset),.i1(intermediate_reg_1[11]),.i2(intermediate_reg_1[10]),.o(intermediate_reg_2[5])); 
fsm fsm_inst_2_895(.clk(clk),.reset(reset),.i1(intermediate_reg_1[9]),.i2(intermediate_reg_1[8]),.o(intermediate_reg_2[4])); 
mux_module mux_module_inst_2_896(.clk(clk),.reset(reset),.i1(intermediate_reg_1[7]),.i2(intermediate_reg_1[6]),.o(intermediate_reg_2[3]),.sel(intermediate_reg_1[0])); 
fsm fsm_inst_2_897(.clk(clk),.reset(reset),.i1(intermediate_reg_1[5]),.i2(intermediate_reg_1[4]),.o(intermediate_reg_2[2])); 
fsm fsm_inst_2_898(.clk(clk),.reset(reset),.i1(intermediate_reg_1[3]),.i2(intermediate_reg_1[2]),.o(intermediate_reg_2[1])); 
mux_module mux_module_inst_2_899(.clk(clk),.reset(reset),.i1(intermediate_reg_1[1]),.i2(intermediate_reg_1[0]),.o(intermediate_reg_2[0]),.sel(intermediate_reg_1[0])); 
always@(posedge clk) begin 
outp [899:0] <= intermediate_reg_2; 
outp[1547:900] <= intermediate_reg_2[647:0] ; 
end 
endmodule 
 

module dpram_2048_40bit_module_4(input clk, input reset, input[415:0] inp, output reg [319:0] outp); 

dpram_2048_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[103:0]),.outp(outp[79:0])); 

dpram_2048_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[207:104]),.outp(outp[159:80])); 

dpram_2048_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[311:208]),.outp(outp[239:160])); 

dpram_2048_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[415:312]),.outp(outp[319:240])); 

endmodule 

module dsp_chain_4_fp16_sop2_mult_module_8(input clk, input reset, input[2047:0] inp, output reg [255:0] outp); 

dsp_chain_4_fp16_sop2_mult_module inst_0 (.clk(clk),.reset(reset),.inp(inp[255:0]),.outp(outp[31:0])); 

dsp_chain_4_fp16_sop2_mult_module inst_1 (.clk(clk),.reset(reset),.inp(inp[511:256]),.outp(outp[63:32])); 

dsp_chain_4_fp16_sop2_mult_module inst_2 (.clk(clk),.reset(reset),.inp(inp[767:512]),.outp(outp[95:64])); 

dsp_chain_4_fp16_sop2_mult_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1023:768]),.outp(outp[127:96])); 

dsp_chain_4_fp16_sop2_mult_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1279:1024]),.outp(outp[159:128])); 

dsp_chain_4_fp16_sop2_mult_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1535:1280]),.outp(outp[191:160])); 

dsp_chain_4_fp16_sop2_mult_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1791:1536]),.outp(outp[223:192])); 

dsp_chain_4_fp16_sop2_mult_module inst_7 (.clk(clk),.reset(reset),.inp(inp[2047:1792]),.outp(outp[255:224])); 

endmodule 

module dsp_chain_2_fp16_sop2_mult_module_4(input clk, input reset, input[511:0] inp, output reg [127:0] outp); 

dsp_chain_2_fp16_sop2_mult_module inst_0 (.clk(clk),.reset(reset),.inp(inp[127:0]),.outp(outp[31:0])); 

dsp_chain_2_fp16_sop2_mult_module inst_1 (.clk(clk),.reset(reset),.inp(inp[255:128]),.outp(outp[63:32])); 

dsp_chain_2_fp16_sop2_mult_module inst_2 (.clk(clk),.reset(reset),.inp(inp[383:256]),.outp(outp[95:64])); 

dsp_chain_2_fp16_sop2_mult_module inst_3 (.clk(clk),.reset(reset),.inp(inp[511:384]),.outp(outp[127:96])); 

endmodule 

module dsp_chain_3_fp16_sop2_mult_module_6(input clk, input reset, input[1151:0] inp, output reg [191:0] outp); 

dsp_chain_3_fp16_sop2_mult_module inst_0 (.clk(clk),.reset(reset),.inp(inp[191:0]),.outp(outp[31:0])); 

dsp_chain_3_fp16_sop2_mult_module inst_1 (.clk(clk),.reset(reset),.inp(inp[383:192]),.outp(outp[63:32])); 

dsp_chain_3_fp16_sop2_mult_module inst_2 (.clk(clk),.reset(reset),.inp(inp[575:384]),.outp(outp[95:64])); 

dsp_chain_3_fp16_sop2_mult_module inst_3 (.clk(clk),.reset(reset),.inp(inp[767:576]),.outp(outp[127:96])); 

dsp_chain_3_fp16_sop2_mult_module inst_4 (.clk(clk),.reset(reset),.inp(inp[959:768]),.outp(outp[159:128])); 

dsp_chain_3_fp16_sop2_mult_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1151:960]),.outp(outp[191:160])); 

endmodule 

module activation_32_8bit_module_4(input clk, input reset, input[1043:0] inp, output reg [1031:0] outp); 

activation_32_8bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[260:0]),.outp(outp[257:0])); 

activation_32_8bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[521:261]),.outp(outp[515:258])); 

activation_32_8bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[782:522]),.outp(outp[773:516])); 

activation_32_8bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1043:783]),.outp(outp[1031:774])); 

endmodule 

module activation_32_16bit_module_3(input clk, input reset, input[1547:0] inp, output reg [1541:0] outp); 

activation_32_16bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[515:0]),.outp(outp[513:0])); 

activation_32_16bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[1031:516]),.outp(outp[1027:514])); 

activation_32_16bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[1547:1032]),.outp(outp[1541:1028])); 

endmodule 

module tanh_16bit_12(input clk, input reset, input[191:0] inp, output reg [191:0] outp); 

tanh_16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[15:0]),.outp(outp[15:0])); 

tanh_16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[31:16]),.outp(outp[31:16])); 

tanh_16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[47:32]),.outp(outp[47:32])); 

tanh_16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[63:48]),.outp(outp[63:48])); 

tanh_16bit inst_4 (.clk(clk),.reset(reset),.inp(inp[79:64]),.outp(outp[79:64])); 

tanh_16bit inst_5 (.clk(clk),.reset(reset),.inp(inp[95:80]),.outp(outp[95:80])); 

tanh_16bit inst_6 (.clk(clk),.reset(reset),.inp(inp[111:96]),.outp(outp[111:96])); 

tanh_16bit inst_7 (.clk(clk),.reset(reset),.inp(inp[127:112]),.outp(outp[127:112])); 

tanh_16bit inst_8 (.clk(clk),.reset(reset),.inp(inp[143:128]),.outp(outp[143:128])); 

tanh_16bit inst_9 (.clk(clk),.reset(reset),.inp(inp[159:144]),.outp(outp[159:144])); 

tanh_16bit inst_10 (.clk(clk),.reset(reset),.inp(inp[175:160]),.outp(outp[175:160])); 

tanh_16bit inst_11 (.clk(clk),.reset(reset),.inp(inp[191:176]),.outp(outp[191:176])); 

endmodule 

module activation_32_8bit_module_6(input clk, input reset, input[1565:0] inp, output reg [1547:0] outp); 

activation_32_8bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[260:0]),.outp(outp[257:0])); 

activation_32_8bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[521:261]),.outp(outp[515:258])); 

activation_32_8bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[782:522]),.outp(outp[773:516])); 

activation_32_8bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1043:783]),.outp(outp[1031:774])); 

activation_32_8bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1304:1044]),.outp(outp[1289:1032])); 

activation_32_8bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1565:1305]),.outp(outp[1547:1290])); 

endmodule 

module sigmoid_16bit_24(input clk, input reset, input[383:0] inp, output reg [383:0] outp); 

sigmoid_16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[15:0]),.outp(outp[15:0])); 

sigmoid_16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[31:16]),.outp(outp[31:16])); 

sigmoid_16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[47:32]),.outp(outp[47:32])); 

sigmoid_16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[63:48]),.outp(outp[63:48])); 

sigmoid_16bit inst_4 (.clk(clk),.reset(reset),.inp(inp[79:64]),.outp(outp[79:64])); 

sigmoid_16bit inst_5 (.clk(clk),.reset(reset),.inp(inp[95:80]),.outp(outp[95:80])); 

sigmoid_16bit inst_6 (.clk(clk),.reset(reset),.inp(inp[111:96]),.outp(outp[111:96])); 

sigmoid_16bit inst_7 (.clk(clk),.reset(reset),.inp(inp[127:112]),.outp(outp[127:112])); 

sigmoid_16bit inst_8 (.clk(clk),.reset(reset),.inp(inp[143:128]),.outp(outp[143:128])); 

sigmoid_16bit inst_9 (.clk(clk),.reset(reset),.inp(inp[159:144]),.outp(outp[159:144])); 

sigmoid_16bit inst_10 (.clk(clk),.reset(reset),.inp(inp[175:160]),.outp(outp[175:160])); 

sigmoid_16bit inst_11 (.clk(clk),.reset(reset),.inp(inp[191:176]),.outp(outp[191:176])); 

sigmoid_16bit inst_12 (.clk(clk),.reset(reset),.inp(inp[207:192]),.outp(outp[207:192])); 

sigmoid_16bit inst_13 (.clk(clk),.reset(reset),.inp(inp[223:208]),.outp(outp[223:208])); 

sigmoid_16bit inst_14 (.clk(clk),.reset(reset),.inp(inp[239:224]),.outp(outp[239:224])); 

sigmoid_16bit inst_15 (.clk(clk),.reset(reset),.inp(inp[255:240]),.outp(outp[255:240])); 

sigmoid_16bit inst_16 (.clk(clk),.reset(reset),.inp(inp[271:256]),.outp(outp[271:256])); 

sigmoid_16bit inst_17 (.clk(clk),.reset(reset),.inp(inp[287:272]),.outp(outp[287:272])); 

sigmoid_16bit inst_18 (.clk(clk),.reset(reset),.inp(inp[303:288]),.outp(outp[303:288])); 

sigmoid_16bit inst_19 (.clk(clk),.reset(reset),.inp(inp[319:304]),.outp(outp[319:304])); 

sigmoid_16bit inst_20 (.clk(clk),.reset(reset),.inp(inp[335:320]),.outp(outp[335:320])); 

sigmoid_16bit inst_21 (.clk(clk),.reset(reset),.inp(inp[351:336]),.outp(outp[351:336])); 

sigmoid_16bit inst_22 (.clk(clk),.reset(reset),.inp(inp[367:352]),.outp(outp[367:352])); 

sigmoid_16bit inst_23 (.clk(clk),.reset(reset),.inp(inp[383:368]),.outp(outp[383:368])); 

endmodule 

module activation_32_8bit_module_8(input clk, input reset, input[2087:0] inp, output reg [2063:0] outp); 

activation_32_8bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[260:0]),.outp(outp[257:0])); 

activation_32_8bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[521:261]),.outp(outp[515:258])); 

activation_32_8bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[782:522]),.outp(outp[773:516])); 

activation_32_8bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1043:783]),.outp(outp[1031:774])); 

activation_32_8bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1304:1044]),.outp(outp[1289:1032])); 

activation_32_8bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1565:1305]),.outp(outp[1547:1290])); 

activation_32_8bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1826:1566]),.outp(outp[1805:1548])); 

activation_32_8bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[2087:1827]),.outp(outp[2063:1806])); 

endmodule 

module dpram_4096_40bit_module_10(input clk, input reset, input[1059:0] inp, output reg [799:0] outp); 

dpram_4096_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[105:0]),.outp(outp[79:0])); 

dpram_4096_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[211:106]),.outp(outp[159:80])); 

dpram_4096_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[317:212]),.outp(outp[239:160])); 

dpram_4096_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[423:318]),.outp(outp[319:240])); 

dpram_4096_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[529:424]),.outp(outp[399:320])); 

dpram_4096_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[635:530]),.outp(outp[479:400])); 

dpram_4096_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[741:636]),.outp(outp[559:480])); 

dpram_4096_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[847:742]),.outp(outp[639:560])); 

dpram_4096_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[953:848]),.outp(outp[719:640])); 

dpram_4096_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1059:954]),.outp(outp[799:720])); 

endmodule 

module dpram_4096_60bit_module_8(input clk, input reset, input[1167:0] inp, output reg [959:0] outp); 

dpram_4096_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[145:0]),.outp(outp[119:0])); 

dpram_4096_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[291:146]),.outp(outp[239:120])); 

dpram_4096_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[437:292]),.outp(outp[359:240])); 

dpram_4096_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[583:438]),.outp(outp[479:360])); 

dpram_4096_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[729:584]),.outp(outp[599:480])); 

dpram_4096_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[875:730]),.outp(outp[719:600])); 

dpram_4096_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1021:876]),.outp(outp[839:720])); 

dpram_4096_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1167:1022]),.outp(outp[959:840])); 

endmodule 

module dpram_2048_60bit_module_20(input clk, input reset, input[2879:0] inp, output reg [2399:0] outp); 

dpram_2048_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[143:0]),.outp(outp[119:0])); 

dpram_2048_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[287:144]),.outp(outp[239:120])); 

dpram_2048_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[431:288]),.outp(outp[359:240])); 

dpram_2048_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[575:432]),.outp(outp[479:360])); 

dpram_2048_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[719:576]),.outp(outp[599:480])); 

dpram_2048_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[863:720]),.outp(outp[719:600])); 

dpram_2048_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1007:864]),.outp(outp[839:720])); 

dpram_2048_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1151:1008]),.outp(outp[959:840])); 

dpram_2048_60bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[1295:1152]),.outp(outp[1079:960])); 

dpram_2048_60bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1439:1296]),.outp(outp[1199:1080])); 

dpram_2048_60bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[1583:1440]),.outp(outp[1319:1200])); 

dpram_2048_60bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[1727:1584]),.outp(outp[1439:1320])); 

dpram_2048_60bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[1871:1728]),.outp(outp[1559:1440])); 

dpram_2048_60bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[2015:1872]),.outp(outp[1679:1560])); 

dpram_2048_60bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[2159:2016]),.outp(outp[1799:1680])); 

dpram_2048_60bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[2303:2160]),.outp(outp[1919:1800])); 

dpram_2048_60bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[2447:2304]),.outp(outp[2039:1920])); 

dpram_2048_60bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[2591:2448]),.outp(outp[2159:2040])); 

dpram_2048_60bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[2735:2592]),.outp(outp[2279:2160])); 

dpram_2048_60bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[2879:2736]),.outp(outp[2399:2280])); 

endmodule 

module dpram_2048_40bit_module_24(input clk, input reset, input[2495:0] inp, output reg [1919:0] outp); 

dpram_2048_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[103:0]),.outp(outp[79:0])); 

dpram_2048_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[207:104]),.outp(outp[159:80])); 

dpram_2048_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[311:208]),.outp(outp[239:160])); 

dpram_2048_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[415:312]),.outp(outp[319:240])); 

dpram_2048_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[519:416]),.outp(outp[399:320])); 

dpram_2048_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[623:520]),.outp(outp[479:400])); 

dpram_2048_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[727:624]),.outp(outp[559:480])); 

dpram_2048_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[831:728]),.outp(outp[639:560])); 

dpram_2048_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[935:832]),.outp(outp[719:640])); 

dpram_2048_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1039:936]),.outp(outp[799:720])); 

dpram_2048_40bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[1143:1040]),.outp(outp[879:800])); 

dpram_2048_40bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[1247:1144]),.outp(outp[959:880])); 

dpram_2048_40bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[1351:1248]),.outp(outp[1039:960])); 

dpram_2048_40bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[1455:1352]),.outp(outp[1119:1040])); 

dpram_2048_40bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[1559:1456]),.outp(outp[1199:1120])); 

dpram_2048_40bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[1663:1560]),.outp(outp[1279:1200])); 

dpram_2048_40bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[1767:1664]),.outp(outp[1359:1280])); 

dpram_2048_40bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[1871:1768]),.outp(outp[1439:1360])); 

dpram_2048_40bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[1975:1872]),.outp(outp[1519:1440])); 

dpram_2048_40bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[2079:1976]),.outp(outp[1599:1520])); 

dpram_2048_40bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[2183:2080]),.outp(outp[1679:1600])); 

dpram_2048_40bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[2287:2184]),.outp(outp[1759:1680])); 

dpram_2048_40bit_module inst_22 (.clk(clk),.reset(reset),.inp(inp[2391:2288]),.outp(outp[1839:1760])); 

dpram_2048_40bit_module inst_23 (.clk(clk),.reset(reset),.inp(inp[2495:2392]),.outp(outp[1919:1840])); 

endmodule 

module dpram_4096_40bit_module_22(input clk, input reset, input[2331:0] inp, output reg [1759:0] outp); 

dpram_4096_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[105:0]),.outp(outp[79:0])); 

dpram_4096_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[211:106]),.outp(outp[159:80])); 

dpram_4096_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[317:212]),.outp(outp[239:160])); 

dpram_4096_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[423:318]),.outp(outp[319:240])); 

dpram_4096_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[529:424]),.outp(outp[399:320])); 

dpram_4096_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[635:530]),.outp(outp[479:400])); 

dpram_4096_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[741:636]),.outp(outp[559:480])); 

dpram_4096_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[847:742]),.outp(outp[639:560])); 

dpram_4096_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[953:848]),.outp(outp[719:640])); 

dpram_4096_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1059:954]),.outp(outp[799:720])); 

dpram_4096_40bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[1165:1060]),.outp(outp[879:800])); 

dpram_4096_40bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[1271:1166]),.outp(outp[959:880])); 

dpram_4096_40bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[1377:1272]),.outp(outp[1039:960])); 

dpram_4096_40bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[1483:1378]),.outp(outp[1119:1040])); 

dpram_4096_40bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[1589:1484]),.outp(outp[1199:1120])); 

dpram_4096_40bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[1695:1590]),.outp(outp[1279:1200])); 

dpram_4096_40bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[1801:1696]),.outp(outp[1359:1280])); 

dpram_4096_40bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[1907:1802]),.outp(outp[1439:1360])); 

dpram_4096_40bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[2013:1908]),.outp(outp[1519:1440])); 

dpram_4096_40bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[2119:2014]),.outp(outp[1599:1520])); 

dpram_4096_40bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[2225:2120]),.outp(outp[1679:1600])); 

dpram_4096_40bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[2331:2226]),.outp(outp[1759:1680])); 

endmodule 

module dpram_2048_60bit_module_30(input clk, input reset, input[4319:0] inp, output reg [3599:0] outp); 

dpram_2048_60bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[143:0]),.outp(outp[119:0])); 

dpram_2048_60bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[287:144]),.outp(outp[239:120])); 

dpram_2048_60bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[431:288]),.outp(outp[359:240])); 

dpram_2048_60bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[575:432]),.outp(outp[479:360])); 

dpram_2048_60bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[719:576]),.outp(outp[599:480])); 

dpram_2048_60bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[863:720]),.outp(outp[719:600])); 

dpram_2048_60bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1007:864]),.outp(outp[839:720])); 

dpram_2048_60bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1151:1008]),.outp(outp[959:840])); 

dpram_2048_60bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[1295:1152]),.outp(outp[1079:960])); 

dpram_2048_60bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1439:1296]),.outp(outp[1199:1080])); 

dpram_2048_60bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[1583:1440]),.outp(outp[1319:1200])); 

dpram_2048_60bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[1727:1584]),.outp(outp[1439:1320])); 

dpram_2048_60bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[1871:1728]),.outp(outp[1559:1440])); 

dpram_2048_60bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[2015:1872]),.outp(outp[1679:1560])); 

dpram_2048_60bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[2159:2016]),.outp(outp[1799:1680])); 

dpram_2048_60bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[2303:2160]),.outp(outp[1919:1800])); 

dpram_2048_60bit_module inst_16 (.clk(clk),.reset(reset),.inp(inp[2447:2304]),.outp(outp[2039:1920])); 

dpram_2048_60bit_module inst_17 (.clk(clk),.reset(reset),.inp(inp[2591:2448]),.outp(outp[2159:2040])); 

dpram_2048_60bit_module inst_18 (.clk(clk),.reset(reset),.inp(inp[2735:2592]),.outp(outp[2279:2160])); 

dpram_2048_60bit_module inst_19 (.clk(clk),.reset(reset),.inp(inp[2879:2736]),.outp(outp[2399:2280])); 

dpram_2048_60bit_module inst_20 (.clk(clk),.reset(reset),.inp(inp[3023:2880]),.outp(outp[2519:2400])); 

dpram_2048_60bit_module inst_21 (.clk(clk),.reset(reset),.inp(inp[3167:3024]),.outp(outp[2639:2520])); 

dpram_2048_60bit_module inst_22 (.clk(clk),.reset(reset),.inp(inp[3311:3168]),.outp(outp[2759:2640])); 

dpram_2048_60bit_module inst_23 (.clk(clk),.reset(reset),.inp(inp[3455:3312]),.outp(outp[2879:2760])); 

dpram_2048_60bit_module inst_24 (.clk(clk),.reset(reset),.inp(inp[3599:3456]),.outp(outp[2999:2880])); 

dpram_2048_60bit_module inst_25 (.clk(clk),.reset(reset),.inp(inp[3743:3600]),.outp(outp[3119:3000])); 

dpram_2048_60bit_module inst_26 (.clk(clk),.reset(reset),.inp(inp[3887:3744]),.outp(outp[3239:3120])); 

dpram_2048_60bit_module inst_27 (.clk(clk),.reset(reset),.inp(inp[4031:3888]),.outp(outp[3359:3240])); 

dpram_2048_60bit_module inst_28 (.clk(clk),.reset(reset),.inp(inp[4175:4032]),.outp(outp[3479:3360])); 

dpram_2048_60bit_module inst_29 (.clk(clk),.reset(reset),.inp(inp[4319:4176]),.outp(outp[3599:3480])); 

endmodule 

module dsp_chain_2_fp16_sop2_mult_module_1(input clk, input reset, input[127:0] inp, output reg [31:0] outp); 

dsp_chain_2_fp16_sop2_mult_module inst_0 (.clk(clk),.reset(reset),.inp(inp[127:0]),.outp(outp[31:0])); 

endmodule 

module dpram_4096_40bit_module_16(input clk, input reset, input[1695:0] inp, output reg [1279:0] outp); 

dpram_4096_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[105:0]),.outp(outp[79:0])); 

dpram_4096_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[211:106]),.outp(outp[159:80])); 

dpram_4096_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[317:212]),.outp(outp[239:160])); 

dpram_4096_40bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[423:318]),.outp(outp[319:240])); 

dpram_4096_40bit_module inst_4 (.clk(clk),.reset(reset),.inp(inp[529:424]),.outp(outp[399:320])); 

dpram_4096_40bit_module inst_5 (.clk(clk),.reset(reset),.inp(inp[635:530]),.outp(outp[479:400])); 

dpram_4096_40bit_module inst_6 (.clk(clk),.reset(reset),.inp(inp[741:636]),.outp(outp[559:480])); 

dpram_4096_40bit_module inst_7 (.clk(clk),.reset(reset),.inp(inp[847:742]),.outp(outp[639:560])); 

dpram_4096_40bit_module inst_8 (.clk(clk),.reset(reset),.inp(inp[953:848]),.outp(outp[719:640])); 

dpram_4096_40bit_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1059:954]),.outp(outp[799:720])); 

dpram_4096_40bit_module inst_10 (.clk(clk),.reset(reset),.inp(inp[1165:1060]),.outp(outp[879:800])); 

dpram_4096_40bit_module inst_11 (.clk(clk),.reset(reset),.inp(inp[1271:1166]),.outp(outp[959:880])); 

dpram_4096_40bit_module inst_12 (.clk(clk),.reset(reset),.inp(inp[1377:1272]),.outp(outp[1039:960])); 

dpram_4096_40bit_module inst_13 (.clk(clk),.reset(reset),.inp(inp[1483:1378]),.outp(outp[1119:1040])); 

dpram_4096_40bit_module inst_14 (.clk(clk),.reset(reset),.inp(inp[1589:1484]),.outp(outp[1199:1120])); 

dpram_4096_40bit_module inst_15 (.clk(clk),.reset(reset),.inp(inp[1695:1590]),.outp(outp[1279:1200])); 

endmodule 

module dsp_chain_4_fp16_sop2_mult_module_20(input clk, input reset, input[5119:0] inp, output reg [639:0] outp); 

dsp_chain_4_fp16_sop2_mult_module inst_0 (.clk(clk),.reset(reset),.inp(inp[255:0]),.outp(outp[31:0])); 

dsp_chain_4_fp16_sop2_mult_module inst_1 (.clk(clk),.reset(reset),.inp(inp[511:256]),.outp(outp[63:32])); 

dsp_chain_4_fp16_sop2_mult_module inst_2 (.clk(clk),.reset(reset),.inp(inp[767:512]),.outp(outp[95:64])); 

dsp_chain_4_fp16_sop2_mult_module inst_3 (.clk(clk),.reset(reset),.inp(inp[1023:768]),.outp(outp[127:96])); 

dsp_chain_4_fp16_sop2_mult_module inst_4 (.clk(clk),.reset(reset),.inp(inp[1279:1024]),.outp(outp[159:128])); 

dsp_chain_4_fp16_sop2_mult_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1535:1280]),.outp(outp[191:160])); 

dsp_chain_4_fp16_sop2_mult_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1791:1536]),.outp(outp[223:192])); 

dsp_chain_4_fp16_sop2_mult_module inst_7 (.clk(clk),.reset(reset),.inp(inp[2047:1792]),.outp(outp[255:224])); 

dsp_chain_4_fp16_sop2_mult_module inst_8 (.clk(clk),.reset(reset),.inp(inp[2303:2048]),.outp(outp[287:256])); 

dsp_chain_4_fp16_sop2_mult_module inst_9 (.clk(clk),.reset(reset),.inp(inp[2559:2304]),.outp(outp[319:288])); 

dsp_chain_4_fp16_sop2_mult_module inst_10 (.clk(clk),.reset(reset),.inp(inp[2815:2560]),.outp(outp[351:320])); 

dsp_chain_4_fp16_sop2_mult_module inst_11 (.clk(clk),.reset(reset),.inp(inp[3071:2816]),.outp(outp[383:352])); 

dsp_chain_4_fp16_sop2_mult_module inst_12 (.clk(clk),.reset(reset),.inp(inp[3327:3072]),.outp(outp[415:384])); 

dsp_chain_4_fp16_sop2_mult_module inst_13 (.clk(clk),.reset(reset),.inp(inp[3583:3328]),.outp(outp[447:416])); 

dsp_chain_4_fp16_sop2_mult_module inst_14 (.clk(clk),.reset(reset),.inp(inp[3839:3584]),.outp(outp[479:448])); 

dsp_chain_4_fp16_sop2_mult_module inst_15 (.clk(clk),.reset(reset),.inp(inp[4095:3840]),.outp(outp[511:480])); 

dsp_chain_4_fp16_sop2_mult_module inst_16 (.clk(clk),.reset(reset),.inp(inp[4351:4096]),.outp(outp[543:512])); 

dsp_chain_4_fp16_sop2_mult_module inst_17 (.clk(clk),.reset(reset),.inp(inp[4607:4352]),.outp(outp[575:544])); 

dsp_chain_4_fp16_sop2_mult_module inst_18 (.clk(clk),.reset(reset),.inp(inp[4863:4608]),.outp(outp[607:576])); 

dsp_chain_4_fp16_sop2_mult_module inst_19 (.clk(clk),.reset(reset),.inp(inp[5119:4864]),.outp(outp[639:608])); 

endmodule 

module sigmoid_16bit_30(input clk, input reset, input[479:0] inp, output reg [479:0] outp); 

sigmoid_16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[15:0]),.outp(outp[15:0])); 

sigmoid_16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[31:16]),.outp(outp[31:16])); 

sigmoid_16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[47:32]),.outp(outp[47:32])); 

sigmoid_16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[63:48]),.outp(outp[63:48])); 

sigmoid_16bit inst_4 (.clk(clk),.reset(reset),.inp(inp[79:64]),.outp(outp[79:64])); 

sigmoid_16bit inst_5 (.clk(clk),.reset(reset),.inp(inp[95:80]),.outp(outp[95:80])); 

sigmoid_16bit inst_6 (.clk(clk),.reset(reset),.inp(inp[111:96]),.outp(outp[111:96])); 

sigmoid_16bit inst_7 (.clk(clk),.reset(reset),.inp(inp[127:112]),.outp(outp[127:112])); 

sigmoid_16bit inst_8 (.clk(clk),.reset(reset),.inp(inp[143:128]),.outp(outp[143:128])); 

sigmoid_16bit inst_9 (.clk(clk),.reset(reset),.inp(inp[159:144]),.outp(outp[159:144])); 

sigmoid_16bit inst_10 (.clk(clk),.reset(reset),.inp(inp[175:160]),.outp(outp[175:160])); 

sigmoid_16bit inst_11 (.clk(clk),.reset(reset),.inp(inp[191:176]),.outp(outp[191:176])); 

sigmoid_16bit inst_12 (.clk(clk),.reset(reset),.inp(inp[207:192]),.outp(outp[207:192])); 

sigmoid_16bit inst_13 (.clk(clk),.reset(reset),.inp(inp[223:208]),.outp(outp[223:208])); 

sigmoid_16bit inst_14 (.clk(clk),.reset(reset),.inp(inp[239:224]),.outp(outp[239:224])); 

sigmoid_16bit inst_15 (.clk(clk),.reset(reset),.inp(inp[255:240]),.outp(outp[255:240])); 

sigmoid_16bit inst_16 (.clk(clk),.reset(reset),.inp(inp[271:256]),.outp(outp[271:256])); 

sigmoid_16bit inst_17 (.clk(clk),.reset(reset),.inp(inp[287:272]),.outp(outp[287:272])); 

sigmoid_16bit inst_18 (.clk(clk),.reset(reset),.inp(inp[303:288]),.outp(outp[303:288])); 

sigmoid_16bit inst_19 (.clk(clk),.reset(reset),.inp(inp[319:304]),.outp(outp[319:304])); 

sigmoid_16bit inst_20 (.clk(clk),.reset(reset),.inp(inp[335:320]),.outp(outp[335:320])); 

sigmoid_16bit inst_21 (.clk(clk),.reset(reset),.inp(inp[351:336]),.outp(outp[351:336])); 

sigmoid_16bit inst_22 (.clk(clk),.reset(reset),.inp(inp[367:352]),.outp(outp[367:352])); 

sigmoid_16bit inst_23 (.clk(clk),.reset(reset),.inp(inp[383:368]),.outp(outp[383:368])); 

sigmoid_16bit inst_24 (.clk(clk),.reset(reset),.inp(inp[399:384]),.outp(outp[399:384])); 

sigmoid_16bit inst_25 (.clk(clk),.reset(reset),.inp(inp[415:400]),.outp(outp[415:400])); 

sigmoid_16bit inst_26 (.clk(clk),.reset(reset),.inp(inp[431:416]),.outp(outp[431:416])); 

sigmoid_16bit inst_27 (.clk(clk),.reset(reset),.inp(inp[447:432]),.outp(outp[447:432])); 

sigmoid_16bit inst_28 (.clk(clk),.reset(reset),.inp(inp[463:448]),.outp(outp[463:448])); 

sigmoid_16bit inst_29 (.clk(clk),.reset(reset),.inp(inp[479:464]),.outp(outp[479:464])); 

endmodule 

module dsp_chain_3_fp16_sop2_mult_module_26(input clk, input reset, input[4991:0] inp, output reg [831:0] outp); 

dsp_chain_3_fp16_sop2_mult_module inst_0 (.clk(clk),.reset(reset),.inp(inp[191:0]),.outp(outp[31:0])); 

dsp_chain_3_fp16_sop2_mult_module inst_1 (.clk(clk),.reset(reset),.inp(inp[383:192]),.outp(outp[63:32])); 

dsp_chain_3_fp16_sop2_mult_module inst_2 (.clk(clk),.reset(reset),.inp(inp[575:384]),.outp(outp[95:64])); 

dsp_chain_3_fp16_sop2_mult_module inst_3 (.clk(clk),.reset(reset),.inp(inp[767:576]),.outp(outp[127:96])); 

dsp_chain_3_fp16_sop2_mult_module inst_4 (.clk(clk),.reset(reset),.inp(inp[959:768]),.outp(outp[159:128])); 

dsp_chain_3_fp16_sop2_mult_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1151:960]),.outp(outp[191:160])); 

dsp_chain_3_fp16_sop2_mult_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1343:1152]),.outp(outp[223:192])); 

dsp_chain_3_fp16_sop2_mult_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1535:1344]),.outp(outp[255:224])); 

dsp_chain_3_fp16_sop2_mult_module inst_8 (.clk(clk),.reset(reset),.inp(inp[1727:1536]),.outp(outp[287:256])); 

dsp_chain_3_fp16_sop2_mult_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1919:1728]),.outp(outp[319:288])); 

dsp_chain_3_fp16_sop2_mult_module inst_10 (.clk(clk),.reset(reset),.inp(inp[2111:1920]),.outp(outp[351:320])); 

dsp_chain_3_fp16_sop2_mult_module inst_11 (.clk(clk),.reset(reset),.inp(inp[2303:2112]),.outp(outp[383:352])); 

dsp_chain_3_fp16_sop2_mult_module inst_12 (.clk(clk),.reset(reset),.inp(inp[2495:2304]),.outp(outp[415:384])); 

dsp_chain_3_fp16_sop2_mult_module inst_13 (.clk(clk),.reset(reset),.inp(inp[2687:2496]),.outp(outp[447:416])); 

dsp_chain_3_fp16_sop2_mult_module inst_14 (.clk(clk),.reset(reset),.inp(inp[2879:2688]),.outp(outp[479:448])); 

dsp_chain_3_fp16_sop2_mult_module inst_15 (.clk(clk),.reset(reset),.inp(inp[3071:2880]),.outp(outp[511:480])); 

dsp_chain_3_fp16_sop2_mult_module inst_16 (.clk(clk),.reset(reset),.inp(inp[3263:3072]),.outp(outp[543:512])); 

dsp_chain_3_fp16_sop2_mult_module inst_17 (.clk(clk),.reset(reset),.inp(inp[3455:3264]),.outp(outp[575:544])); 

dsp_chain_3_fp16_sop2_mult_module inst_18 (.clk(clk),.reset(reset),.inp(inp[3647:3456]),.outp(outp[607:576])); 

dsp_chain_3_fp16_sop2_mult_module inst_19 (.clk(clk),.reset(reset),.inp(inp[3839:3648]),.outp(outp[639:608])); 

dsp_chain_3_fp16_sop2_mult_module inst_20 (.clk(clk),.reset(reset),.inp(inp[4031:3840]),.outp(outp[671:640])); 

dsp_chain_3_fp16_sop2_mult_module inst_21 (.clk(clk),.reset(reset),.inp(inp[4223:4032]),.outp(outp[703:672])); 

dsp_chain_3_fp16_sop2_mult_module inst_22 (.clk(clk),.reset(reset),.inp(inp[4415:4224]),.outp(outp[735:704])); 

dsp_chain_3_fp16_sop2_mult_module inst_23 (.clk(clk),.reset(reset),.inp(inp[4607:4416]),.outp(outp[767:736])); 

dsp_chain_3_fp16_sop2_mult_module inst_24 (.clk(clk),.reset(reset),.inp(inp[4799:4608]),.outp(outp[799:768])); 

dsp_chain_3_fp16_sop2_mult_module inst_25 (.clk(clk),.reset(reset),.inp(inp[4991:4800]),.outp(outp[831:800])); 

endmodule 

module activation_32_16bit_module_4(input clk, input reset, input[2063:0] inp, output reg [2055:0] outp); 

activation_32_16bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[515:0]),.outp(outp[513:0])); 

activation_32_16bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[1031:516]),.outp(outp[1027:514])); 

activation_32_16bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[1547:1032]),.outp(outp[1541:1028])); 

activation_32_16bit_module inst_3 (.clk(clk),.reset(reset),.inp(inp[2063:1548]),.outp(outp[2055:1542])); 

endmodule 

module dpram_2048_40bit_module_3(input clk, input reset, input[311:0] inp, output reg [239:0] outp); 

dpram_2048_40bit_module inst_0 (.clk(clk),.reset(reset),.inp(inp[103:0]),.outp(outp[79:0])); 

dpram_2048_40bit_module inst_1 (.clk(clk),.reset(reset),.inp(inp[207:104]),.outp(outp[159:80])); 

dpram_2048_40bit_module inst_2 (.clk(clk),.reset(reset),.inp(inp[311:208]),.outp(outp[239:160])); 

endmodule 

module dsp_chain_3_fp16_sop2_mult_module_50(input clk, input reset, input[9599:0] inp, output reg [1599:0] outp); 

dsp_chain_3_fp16_sop2_mult_module inst_0 (.clk(clk),.reset(reset),.inp(inp[191:0]),.outp(outp[31:0])); 

dsp_chain_3_fp16_sop2_mult_module inst_1 (.clk(clk),.reset(reset),.inp(inp[383:192]),.outp(outp[63:32])); 

dsp_chain_3_fp16_sop2_mult_module inst_2 (.clk(clk),.reset(reset),.inp(inp[575:384]),.outp(outp[95:64])); 

dsp_chain_3_fp16_sop2_mult_module inst_3 (.clk(clk),.reset(reset),.inp(inp[767:576]),.outp(outp[127:96])); 

dsp_chain_3_fp16_sop2_mult_module inst_4 (.clk(clk),.reset(reset),.inp(inp[959:768]),.outp(outp[159:128])); 

dsp_chain_3_fp16_sop2_mult_module inst_5 (.clk(clk),.reset(reset),.inp(inp[1151:960]),.outp(outp[191:160])); 

dsp_chain_3_fp16_sop2_mult_module inst_6 (.clk(clk),.reset(reset),.inp(inp[1343:1152]),.outp(outp[223:192])); 

dsp_chain_3_fp16_sop2_mult_module inst_7 (.clk(clk),.reset(reset),.inp(inp[1535:1344]),.outp(outp[255:224])); 

dsp_chain_3_fp16_sop2_mult_module inst_8 (.clk(clk),.reset(reset),.inp(inp[1727:1536]),.outp(outp[287:256])); 

dsp_chain_3_fp16_sop2_mult_module inst_9 (.clk(clk),.reset(reset),.inp(inp[1919:1728]),.outp(outp[319:288])); 

dsp_chain_3_fp16_sop2_mult_module inst_10 (.clk(clk),.reset(reset),.inp(inp[2111:1920]),.outp(outp[351:320])); 

dsp_chain_3_fp16_sop2_mult_module inst_11 (.clk(clk),.reset(reset),.inp(inp[2303:2112]),.outp(outp[383:352])); 

dsp_chain_3_fp16_sop2_mult_module inst_12 (.clk(clk),.reset(reset),.inp(inp[2495:2304]),.outp(outp[415:384])); 

dsp_chain_3_fp16_sop2_mult_module inst_13 (.clk(clk),.reset(reset),.inp(inp[2687:2496]),.outp(outp[447:416])); 

dsp_chain_3_fp16_sop2_mult_module inst_14 (.clk(clk),.reset(reset),.inp(inp[2879:2688]),.outp(outp[479:448])); 

dsp_chain_3_fp16_sop2_mult_module inst_15 (.clk(clk),.reset(reset),.inp(inp[3071:2880]),.outp(outp[511:480])); 

dsp_chain_3_fp16_sop2_mult_module inst_16 (.clk(clk),.reset(reset),.inp(inp[3263:3072]),.outp(outp[543:512])); 

dsp_chain_3_fp16_sop2_mult_module inst_17 (.clk(clk),.reset(reset),.inp(inp[3455:3264]),.outp(outp[575:544])); 

dsp_chain_3_fp16_sop2_mult_module inst_18 (.clk(clk),.reset(reset),.inp(inp[3647:3456]),.outp(outp[607:576])); 

dsp_chain_3_fp16_sop2_mult_module inst_19 (.clk(clk),.reset(reset),.inp(inp[3839:3648]),.outp(outp[639:608])); 

dsp_chain_3_fp16_sop2_mult_module inst_20 (.clk(clk),.reset(reset),.inp(inp[4031:3840]),.outp(outp[671:640])); 

dsp_chain_3_fp16_sop2_mult_module inst_21 (.clk(clk),.reset(reset),.inp(inp[4223:4032]),.outp(outp[703:672])); 

dsp_chain_3_fp16_sop2_mult_module inst_22 (.clk(clk),.reset(reset),.inp(inp[4415:4224]),.outp(outp[735:704])); 

dsp_chain_3_fp16_sop2_mult_module inst_23 (.clk(clk),.reset(reset),.inp(inp[4607:4416]),.outp(outp[767:736])); 

dsp_chain_3_fp16_sop2_mult_module inst_24 (.clk(clk),.reset(reset),.inp(inp[4799:4608]),.outp(outp[799:768])); 

dsp_chain_3_fp16_sop2_mult_module inst_25 (.clk(clk),.reset(reset),.inp(inp[4991:4800]),.outp(outp[831:800])); 

dsp_chain_3_fp16_sop2_mult_module inst_26 (.clk(clk),.reset(reset),.inp(inp[5183:4992]),.outp(outp[863:832])); 

dsp_chain_3_fp16_sop2_mult_module inst_27 (.clk(clk),.reset(reset),.inp(inp[5375:5184]),.outp(outp[895:864])); 

dsp_chain_3_fp16_sop2_mult_module inst_28 (.clk(clk),.reset(reset),.inp(inp[5567:5376]),.outp(outp[927:896])); 

dsp_chain_3_fp16_sop2_mult_module inst_29 (.clk(clk),.reset(reset),.inp(inp[5759:5568]),.outp(outp[959:928])); 

dsp_chain_3_fp16_sop2_mult_module inst_30 (.clk(clk),.reset(reset),.inp(inp[5951:5760]),.outp(outp[991:960])); 

dsp_chain_3_fp16_sop2_mult_module inst_31 (.clk(clk),.reset(reset),.inp(inp[6143:5952]),.outp(outp[1023:992])); 

dsp_chain_3_fp16_sop2_mult_module inst_32 (.clk(clk),.reset(reset),.inp(inp[6335:6144]),.outp(outp[1055:1024])); 

dsp_chain_3_fp16_sop2_mult_module inst_33 (.clk(clk),.reset(reset),.inp(inp[6527:6336]),.outp(outp[1087:1056])); 

dsp_chain_3_fp16_sop2_mult_module inst_34 (.clk(clk),.reset(reset),.inp(inp[6719:6528]),.outp(outp[1119:1088])); 

dsp_chain_3_fp16_sop2_mult_module inst_35 (.clk(clk),.reset(reset),.inp(inp[6911:6720]),.outp(outp[1151:1120])); 

dsp_chain_3_fp16_sop2_mult_module inst_36 (.clk(clk),.reset(reset),.inp(inp[7103:6912]),.outp(outp[1183:1152])); 

dsp_chain_3_fp16_sop2_mult_module inst_37 (.clk(clk),.reset(reset),.inp(inp[7295:7104]),.outp(outp[1215:1184])); 

dsp_chain_3_fp16_sop2_mult_module inst_38 (.clk(clk),.reset(reset),.inp(inp[7487:7296]),.outp(outp[1247:1216])); 

dsp_chain_3_fp16_sop2_mult_module inst_39 (.clk(clk),.reset(reset),.inp(inp[7679:7488]),.outp(outp[1279:1248])); 

dsp_chain_3_fp16_sop2_mult_module inst_40 (.clk(clk),.reset(reset),.inp(inp[7871:7680]),.outp(outp[1311:1280])); 

dsp_chain_3_fp16_sop2_mult_module inst_41 (.clk(clk),.reset(reset),.inp(inp[8063:7872]),.outp(outp[1343:1312])); 

dsp_chain_3_fp16_sop2_mult_module inst_42 (.clk(clk),.reset(reset),.inp(inp[8255:8064]),.outp(outp[1375:1344])); 

dsp_chain_3_fp16_sop2_mult_module inst_43 (.clk(clk),.reset(reset),.inp(inp[8447:8256]),.outp(outp[1407:1376])); 

dsp_chain_3_fp16_sop2_mult_module inst_44 (.clk(clk),.reset(reset),.inp(inp[8639:8448]),.outp(outp[1439:1408])); 

dsp_chain_3_fp16_sop2_mult_module inst_45 (.clk(clk),.reset(reset),.inp(inp[8831:8640]),.outp(outp[1471:1440])); 

dsp_chain_3_fp16_sop2_mult_module inst_46 (.clk(clk),.reset(reset),.inp(inp[9023:8832]),.outp(outp[1503:1472])); 

dsp_chain_3_fp16_sop2_mult_module inst_47 (.clk(clk),.reset(reset),.inp(inp[9215:9024]),.outp(outp[1535:1504])); 

dsp_chain_3_fp16_sop2_mult_module inst_48 (.clk(clk),.reset(reset),.inp(inp[9407:9216]),.outp(outp[1567:1536])); 

dsp_chain_3_fp16_sop2_mult_module inst_49 (.clk(clk),.reset(reset),.inp(inp[9599:9408]),.outp(outp[1599:1568])); 

endmodule 


module adder_tree_3_fp16bit_4(input clk, input reset, input[527:0] inp, output reg [63:0] outp); 

adder_tree_3_fp16bit inst_0 (.clk(clk),.reset(reset),.inp(inp[131:0]),.outp(outp[15:0])); 

adder_tree_3_fp16bit inst_1 (.clk(clk),.reset(reset),.inp(inp[263:132]),.outp(outp[31:16])); 

adder_tree_3_fp16bit inst_2 (.clk(clk),.reset(reset),.inp(inp[395:264]),.outp(outp[47:32])); 

adder_tree_3_fp16bit inst_3 (.clk(clk),.reset(reset),.inp(inp[527:396]),.outp(outp[63:48])); 

endmodule 


module adder_tree_1_16bit (input clk,input reset,input [31:0] inp, output reg [31:0] outp);

adder_tree_1stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.sum_out(outp));

endmodule

module adder_tree_2_16bit (input clk, input reset, input [63:0] inp, output reg [31:0] outp);

adder_tree_2stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.sum_out(outp));

endmodule

module adder_tree_3_16bit (input clk, input reset, input [127:0] inp, output reg [31:0] outp);

adder_tree_3stage_16bit inst (.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.inp20(inp[79:64]),.inp21(inp[95:80]),.inp30(inp[111:96]),.inp31(inp[127:112]),.sum_out(outp));

endmodule

module adder_tree_4_16bit (input clk, input reset, input [255:0] inp, output reg [31:0] outp);

adder_tree_4stage_16bit inst(.clk(clk),.reset(reset),.inp00(inp[15:0]),.inp01(inp[31:16]),.inp10(inp[47:32]),.inp11(inp[63:48]),.inp20(inp[79:64]),.inp21(inp[95:80]),.inp30(inp[111:96]),.inp31(inp[127:112]),.inp40(inp[143:128]),.inp41(inp[159:144]),.inp50(inp[175:160]),.inp51(inp[191:176]),.inp60(inp[207:192]),.inp61(inp[223:208]),.inp70(inp[239:224]),.inp71(inp[255:240]),.sum_out(outp));

endmodule

module adder_tree_1_8bit (input clk, input reset, input [15:0] inp, output reg [15:0] outp);

adder_tree_1stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.sum_out(outp));

endmodule

module adder_tree_2_8bit (input clk, input reset, input [31:0] inp, output reg [15:0] outp);

adder_tree_2stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.sum_out(outp));

endmodule

module adder_tree_3_8bit (input clk, input reset, input [63:0] inp, output reg [15:0] outp);

adder_tree_3stage_8bit inst (.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.inp20(inp[39:32]),.inp21(inp[47:40]),.inp30(inp[55:48]),.inp31(inp[63:56]),.sum_out(outp));

endmodule

module adder_tree_4_8bit (input clk, input reset, input [127:0] inp, output reg [15:0] outp);

adder_tree_4stage_8bit inst(.clk(clk),.reset(reset),.inp00(inp[7:0]),.inp01(inp[15:8]),.inp10(inp[23:16]),.inp11(inp[31:24]),.inp20(inp[39:32]),.inp21(inp[47:40]),.inp30(inp[55:48]),.inp31(inp[63:56]),.inp40(inp[71:64]),.inp41(inp[79:72]),.inp50(inp[87:80]),.inp51(inp[95:88]),.inp60(inp[103:96]),.inp61(inp[111:104]),.inp70(inp[119:112]),.inp71(inp[127:120]),.sum_out(outp));

endmodule

module adder_tree_1_4bit (input clk, input reset, input [7:0] inp, output reg [7:0] outp);

adder_tree_1stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.sum_out(outp));

endmodule

module adder_tree_2_4bit (input clk, input reset, input [15:0] inp, output reg [7:0] outp);

adder_tree_2stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.sum_out(outp));

endmodule

module adder_tree_3_4bit (input clk, input reset, input [31:0] inp, output reg [7:0] outp);

adder_tree_3stage_4bit inst (.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.inp20(inp[19:16]),.inp21(inp[23:20]),.inp30(inp[27:24]),.inp31(inp[31:28]),.sum_out(outp));

endmodule

module adder_tree_4_4bit (input clk, input reset, input [63:0] inp, output reg [7:0] outp);

adder_tree_4stage_4bit inst(.clk(clk),.reset(reset),.inp00(inp[3:0]),.inp01(inp[7:4]),.inp10(inp[11:8]),.inp11(inp[15:12]),.inp20(inp[19:16]),.inp21(inp[23:20]),.inp30(inp[27:24]),.inp31(inp[31:28]),.inp40(inp[35:32]),.inp41(inp[39:36]),.inp50(inp[43:40]),.inp51(inp[47:44]),.inp60(inp[51:48]),.inp61(inp[55:52]),.inp70(inp[59:56]),.inp71(inp[63:60]),.sum_out(outp));

endmodule

module adder_tree_3_fp16bit (input clk, input reset, input [131:0] inp, output reg [15:0] outp);

mode4_adder_tree inst(
  .inp0(inp[15:0]),
  .inp1(inp[31:16]),
  .inp2(inp[47:32]),
  .inp3(inp[63:48]),
  .inp4(inp[79:64]),
  .inp5(inp[95:80]),
  .inp6(inp[111:96]),
  .inp7(inp[127:112]),
  .mode4_stage0_run(inp[128]),
  .mode4_stage1_run(inp[129]),
  .mode4_stage2_run(inp[130]),
  .mode4_stage3_run(inp[131]),

  .clk(clk),
  .reset(reset),
  .outp(outp[15:0])
);

endmodule

module dpram_1024_32bit_module (input clk, input reset, input [85:0] inp, output reg [63:0] outp);

dpram inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[53:22]),.data_b(inp[85:54]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_1024_64bit_module (input clk, input reset, input [149:0] inp, output reg [63:0] outp );

dpram_1024_64bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[85:22]),.data_b(inp[149:86]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_2048_64bit_module (input clk, input reset, input [151:0] inp, output reg [127:0] outp);

dpram_2048_64bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[87:24]),.data_b(inp[151:88]),.out_a(outp[63:0]),.out_b(outp[127:64]));

endmodule

module dpram_2048_32bit_module (input clk, input reset, input [87:0] inp, output reg [63:0] outp);

dpram_2048_32bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[55:24]),.data_b(inp[87:56]),.out_a(outp[31:0]),.out_b(outp[63:32]));

endmodule

module dpram_1024_40bit_module (input clk, input reset, input [101:0] inp, output reg [79:0] outp);

dpram_1024_40bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[61:22]),.data_b(inp[101:62]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_1024_60bit_module (input clk, input reset, input [141:0] inp, output reg [119:0] outp);

dpram_1024_60bit inst (.clk(clk),.address_a(inp[9:0]),.address_b(inp[19:10]),.wren_a(inp[20]),.wren_b(inp[21]),.data_a(inp[81:22]),.data_b(inp[141:82]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dpram_2048_40bit_module (input clk, input reset, input [103:0] inp, output reg [79:0] outp);

dpram_2048_40bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[63:24]),.data_b(inp[103:64]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_2048_60bit_module (input clk, input reset, input [143:0] inp, output reg [119:0] outp);

dpram_2048_60bit inst (.clk(clk),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[83:24]),.data_b(inp[143:84]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dpram_4096_40bit_module (input clk, input reset, input [105:0] inp, output reg [79:0] outp);

dpram_4096_40bit inst (.clk(clk),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[65:26]),.data_b(inp[105:66]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dpram_4096_60bit_module (input clk, input reset, input [145:0] inp, output reg [119:0] outp);

dpram_4096_60bit inst (.clk(clk),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[85:26]),.data_b(inp[145:86]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module spram_1024_32bit_module (input clk,input reset,input [42:0] inp, output reg [31:0] outp);

spram inst (.clk(clk),.address(inp[9:0]),.wren(inp[10]),.data(inp[42:11]),.out(outp));

endmodule

module spram_2048_40bit_module (input clk,input reset,input [51:0] inp, output reg [39:0] outp);

spram_2048_40bit inst (.clk(clk),.address(inp[10:0]),.wren(inp[11]),.data(inp[51:12]),.out(outp));

endmodule

module spram_2048_60bit_module (input clk,input reset,input [71:0] inp, output reg [59:0] outp);

spram_2048_60bit inst (.clk(clk),.address(inp[10:0]),.wren(inp[11]),.data(inp[71:12]),.out(outp));

endmodule

module spram_4096_40bit_module (input clk,input reset,input [52:0] inp, output reg [39:0] outp);

spram_4096_40bit inst (.clk(clk),.address(inp[11:0]),.wren(inp[12]),.data(inp[52:13]),.out(outp));

endmodule

module spram_4096_60bit_module (input clk,input reset,input [72:0] inp, output reg [59:0] outp);

spram_4096_60bit inst (.clk(clk),.address(inp[11:0]),.wren(inp[12]),.data(inp[72:13]),.out(outp));

endmodule

module dbram_2048_40bit_module (input clk,input reset,input [103:0] inp, output reg [79:0] outp);

dbram_2048_40bit inst (.clk(clk),.reset(reset),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[63:24]),.data_b(inp[103:64]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dbram_2048_60bit_module (input clk,input reset,input [143:0] inp, output reg [119:0] outp);

dbram_2048_60bit inst (.clk(clk),.reset(reset),.address_a(inp[10:0]),.address_b(inp[21:11]),.wren_a(inp[22]),.wren_b(inp[23]),.data_a(inp[83:24]),.data_b(inp[143:84]),.out_a(outp[59:0]),.out_b(outp[119:60]));

endmodule

module dbram_4096_40bit_module (input clk,input reset,input [105:0] inp, output reg [79:0] outp);

dbram_4096_40bit inst (.clk(clk),.reset(reset),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[65:26]),.data_b(inp[105:66]),.out_a(outp[39:0]),.out_b(outp[79:40]));

endmodule

module dbram_4096_60bit_module (input clk,input reset,input [145:0] inp, output reg [119:0] outp);

dbram_4096_60bit inst (.clk(clk),.reset(reset),.address_a(inp[11:0]),.address_b(inp[23:12]),.wren_a(inp[24]),.wren_b(inp[25]),.data_a(inp[85:26]),.data_b(inp[145:86]),.out_a(outp[59:0]),.out_b(outp[119:40]));

endmodule


module fifo_256_40bit_module (input clk,input reset,input [42:0] inp, output reg [41:0] outp);

fifo_256_40bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[40:1]),.we(inp[41]),.dout(outp[39:0]),.re(inp[42]),.full(outp[40]),.empty(outp[41]));

endmodule

module fifo_256_60bit_module (input clk,input reset,input [62:0] inp, output reg [61:0] outp);

fifo_256_60bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[60:1]),.we(inp[61]),.dout(outp[59:0]),.re(inp[62]),.full(outp[60]),.empty(outp[61]));

endmodule

module fifo_512_60bit_module (input clk,input reset,input [62:0] inp, output reg [61:0] outp);

fifo_512_60bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[60:1]),.we(inp[61]),.dout(outp[59:0]),.re(inp[62]),.full(outp[60]),.empty(outp[61]));

endmodule

module fifo_512_40bit_module (input clk,input reset,input [42:0] inp, output reg [41:0] outp);

fifo_512_40bit inst (.clk(clk),.rst(reset),.clr(inp[0]),.din(inp[40:1]),.we(inp[41]),.dout(outp[39:0]),.re(inp[42]),.full(outp[40]),.empty(outp[41]));

endmodule

module tanh_16bit (input clk,input reset, input [15:0] inp, output reg [15:0] outp);

tanh inst (.x(inp),.tanh_out(outp));

endmodule

module sigmoid_16bit (input clk,input reset, input [15:0] inp, output reg [15:0] outp);

sigmoid inst (.x(inp),.sig_out(outp));

endmodule

module systolic_array_4_16bit (input clk, input reset, input [254:0] inp, output reg [130:0] outp);

matmul_4x4_systolic inst(
 .clk(clk),
 .reset(inp[254]),
 .pe_reset(reset),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[11:1]),
 .address_mat_b(inp[22:12]),
 .address_mat_c(inp[33:23]),
 .address_stride_a(inp[41:34]),
 .address_stride_b(inp[49:42]),
 .address_stride_c(inp[57:50]),
 .a_data(inp[89:58]),
 .b_data(inp[121:90]),
 .a_data_in(inp[153:122]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[185:154]),
 .c_data_in(inp[217:186]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[32:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[64:33]),
 .b_data_out(outp[96:65]),
 .a_addr(outp[107:97]),
 .b_addr(outp[118:108]),
 .c_addr(outp[129:119]),
 .c_data_available(outp[130]),
 .validity_mask_a_rows(inp[221:218]),
 .validity_mask_a_cols_b_rows(inp[225:222]),
 .validity_mask_b_cols(inp[229:226]),
 .final_mat_mul_size(inp[237:230]),
 .a_loc(inp[245:238]),
 .b_loc(inp[253:246])
);

endmodule

module systolic_array_8_16bit (input clk, input reset, input [785:0] inp, output reg [433:0] outp);

matmul_8x8_systolic inst(
 .clk(clk),
 .reset(reset),
 .pe_reset(inp[785]),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[16:1]),
 .address_mat_b(inp[32:17]),
 .address_mat_c(inp[48:33]),
 .address_stride_a(inp[64:49]),
 .address_stride_b(inp[80:65]),
 .address_stride_c(inp[96:81]),
 .a_data(inp[224:97]),
 .b_data(inp[352:225]),
 .a_data_in(inp[480:353]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[608:481]),
 .c_data_in(inp[736:609]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[128:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[256:129]),
 .b_data_out(outp[384:257]),
 .a_addr(outp[400:385]),
 .b_addr(outp[416:401]),
 .c_addr(outp[432:417]),
 .c_data_available(outp[433]),
 .validity_mask_a_rows(inp[744:737]),
 .validity_mask_a_cols_b_rows(inp[752:745]),
 .validity_mask_b_cols(inp[760:753]),
 .final_mat_mul_size(inp[768:761]),
 .a_loc(inp[776:769]),
 .b_loc(inp[784:777])
);

endmodule

module systolic_array_4_fp16bit (input clk, input reset, input [417:0] inp, output reg [223:0] outp);

matmul_4x4_fp_systolic inst(
 .clk(clk),
 .reset(reset),
 .pe_reset(inp[417]),
 .start_mat_mul(inp[0]),
 .done_mat_mul(outp[0]),
 .address_mat_a(inp[10:1]),
 .address_mat_b(inp[20:11]),
 .address_mat_c(inp[30:21]),
 .address_stride_a(inp[40:31]),
 .address_stride_b(inp[50:41]),
 .address_stride_c(inp[60:51]),
 .a_data(inp[124:61]),
 .b_data(inp[188:125]),
 .a_data_in(inp[252:189]), //Data values coming in from previous matmul - systolic connections
 .b_data_in(inp[316:253]),
 .c_data_in(inp[380:317]), //Data values coming in from previous matmul - systolic shifting
 .c_data_out(outp[64:1]), //Data values going out to next matmul - systolic shifting
 .a_data_out(outp[128:65]),
 .b_data_out(outp[192:129]),
 .a_addr(outp[202:193]),
 .b_addr(outp[212:203]),
 .c_addr(outp[222:213]),
 .c_data_available(outp[223]),
 .validity_mask_a_rows(inp[384:381]),
 .validity_mask_a_cols_b_rows(inp[388:385]),
 .validity_mask_b_cols(inp[392:389]),
 .final_mat_mul_size(inp[400:393]),
 .a_loc(inp[408:401]),
 .b_loc(inp[416:409])
);

endmodule

module dsp_chain_2_int_sop_2_module (input clk, input reset, input [147:0] inp, output reg [36:0] outp);

dsp_chain_2_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.result(outp[36:0]));

endmodule

module dsp_chain_3_int_sop_2_module (input clk, input reset, input [221:0] inp, output reg [36:0] outp);

dsp_chain_3_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.ax3(inp[165:148]),.ay3(inp[184:166]),.bx3(inp[202:185]),.by3(inp[221:203]),.result(outp[36:0]));

endmodule

module dsp_chain_4_int_sop_2_module (input clk, input reset, input [295:0] inp, output reg [36:0] outp);

dsp_chain_4_int_sop_2 inst(.clk(clk),.reset(reset),.ax1(inp[17:0]),.ay1(inp[36:18]),.bx1(inp[54:37]),.by1(inp[73:55]),.ax2(inp[91:74]),.ay2(inp[110:92]),.bx2(inp[128:111]),.by2(inp[147:129]),.ax3(inp[165:148]),.ay3(inp[184:166]),.bx3(inp[202:185]),.by3(inp[221:203]),.ax4(inp[239:222]),.ay4(inp[258:240]),.bx4(inp[276:259]),.by4(inp[295:277]),.result(outp[36:0]));

endmodule

module dsp_chain_2_fp16_sop2_mult_module (input clk, input reset, input [127:0] inp, output reg [31:0] outp);

dsp_chain_2_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.result(outp));

endmodule

module dsp_chain_3_fp16_sop2_mult_module (input clk, input reset, input [191:0] inp, output reg [31:0] outp);

dsp_chain_3_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.top_a3(inp[143:128]),.top_b3(inp[159:144]),.bot_a3(inp[175:160]),.bot_b3(inp[191:176]),.result(outp));

endmodule

module dsp_chain_4_fp16_sop2_mult_module (input clk, input reset, input [255:0] inp, output reg [31:0] outp);

dsp_chain_4_fp16_sop2_mult inst(.clk(clk),.reset(reset),.top_a1(inp[15:0]),.top_b1(inp[31:16]),.bot_a1(inp[47:32]),.bot_b1(inp[63:48]),.top_a2(inp[79:64]),.top_b2(inp[95:80]),.bot_a2(inp[111:96]),.bot_b2(inp[127:112]),.top_a3(inp[143:128]),.top_b3(inp[159:144]),.bot_a3(inp[175:160]),.bot_b3(inp[191:176]),.top_a4(inp[207:192]),.top_b4(inp[223:208]),.bot_a4(inp[239:224]),.bot_b4(inp[255:240]),.result(outp));

endmodule

module tensor_block_bf16_module (input clk, input reset, input [264:0] inp, output reg [271:0] outp);

tensor_block_bf16 inst(
	.clk(clk),
	.reset(reset),

	.data_in(inp[79:0]),
	.cascade_in(inp[159:80]),
	.acc0_in(inp[191:160]),
	.acc1_in(inp[223:192]),
	.acc2_in(inp[255:224]),
	.accumulator_input1_select(inp[258:256]),

	.out0(outp[31:0]),
	.out1(outp[63:32]),
	.out2(outp[95:64]),
	.cascade_out(outp[175:96]),
	.acc0_out(outp[207:176]),
	.acc1_out(outp[239:208]),
	.acc2_out(outp[271:240]),

	.mux1_select(inp[259]),
	.dot_unit_input_1_enable(inp[260]),
	.bank0_data_in_enable(inp[261]),
	.bank1_data_in_enable(inp[262]),
	.cascade_out_select(inp[263]),
	.dot_unit_input_2_select(inp[264])

	);

endmodule

module tensor_block_int8_module (input clk, input reset, input [264:0] inp, output reg [250:0] outp);

tensor_block inst(
	.clk(clk),
	.reset(reset),

	.data_in(inp[79:0]),
	.cascade_in(inp[159:80]),
	.acc0_in(inp[191:160]),
	.acc1_in(inp[223:192]),
	.acc2_in(inp[255:224]),
	.accumulator_input1_select(inp[258:256]),

	.out0(outp[24:0]),
	.out1(outp[49:25]),
	.out2(outp[74:50]),
	.cascade_out(outp[154:75]),
	.acc0_out(outp[186:155]),
	.acc1_out(outp[218:187]),
	.acc2_out(outp[250:219]),

	.mux1_select(inp[259]),
	.dot_unit_input_1_enable(inp[260]),
	.bank0_data_in_enable(inp[261]),
	.bank1_data_in_enable(inp[262]),
	.cascade_out_select(inp[263]),
	.dot_unit_input_2_select(inp[264])

	);

endmodule


module activation_32_8bit_module (input clk, input reset, input [260:0] inp, output reg [257:0] outp);

activation_32_8bit inst (
    .activation_type(inp[0]),
    .enable_activation(inp[1]),
    .in_data_available(inp[2]),
    .inp_data(inp[258:3]),
    .out_data(outp[255:0]),
    .out_data_available(outp[256]),
    .validity_mask(inp[260:259]),
    .done_activation(outp[257]),
    .clk(clk),
    .reset(reset)
);

endmodule

module activation_32_16bit_module (input clk, input reset, input [515:0] inp, output reg [513:0] outp);

activation_32_16bit inst (
    .activation_type(inp[0]),
    .enable_activation(inp[1]),
    .in_data_available(inp[2]),
    .inp_data(inp[514:3]),
    .out_data(outp[511:0]),
    .out_data_available(outp[512]),
    .validity_mask(inp[515:514]),
    .done_activation(outp[513]),
    .clk(clk),
    .reset(reset)
);

endmodule

module fsm(input clk, input reset, input i1, input i2, output reg o);
// mealy machine

reg [1:0] current_state; 
reg [1:0] next_state;

wire [1:0] inp; 
assign inp = {i2,i1}; 

always@(posedge clk) begin 
	if (reset == 1'b1) begin 
		current_state <= 1'b0; 
	end
	else begin 
		current_state <= next_state; 
	end
end

always@(posedge clk) begin 

	next_state = current_state; 

	case(current_state)
		2'b00:	begin 
							if(inp == 2'b00) begin 
								next_state <= 2'b00; 
								o <= 1'b0; 
							end
							if (inp == 2'b01) begin 
								next_state <= 2'b11;
								o <= 1'b1;
							end
							if(inp == 2'b10) begin
  							next_state <= 2'b01;
  							o <= 1'b0;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b10;
							  o <= 1'b0;
							end
					 	end 
		2'b01:	begin 
							if(inp == 2'b00) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b01;
							  o <= 1'b0;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b00;
							  o <= 1'b1;
							end
						end
		2'b10:	begin 
							if(inp == 2'b00) begin
							  next_state <= 2'b11;
							  o <= 1'b0;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b11;
							  o <= 1'b0;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
						end
		2'b11:	begin 
							if(inp == 2'b00) begin
  							next_state <= 2'b00;
							  o <= 1'b1;
							end
							if(inp == 2'b01) begin
							  next_state <= 2'b11;
							  o <= 1'b1;
							end
							if(inp == 2'b10) begin
							  next_state <= 2'b10;
							  o <= 1'b1;
							end
							if(inp == 2'b11) begin
							  next_state <= 2'b01;
							  o <= 1'b1;
							end
						end
//		defualt:	begin  
//								next_state <= 2'b00;
//								o <= 1'b0; 
//							end
	endcase
end 

endmodule 
module xor_module (input clk, input reset, input i1, input i2, output reg o);

always@(posedge clk) begin 
if (reset ==1'b1) begin 
o<= 1'b0; 
end
else begin
o <= i1^i2; 
end 
end
endmodule
module mux_module (input clk, input reset, input i1, input i2, output reg o, input sel);

always@(posedge clk) begin 
if (reset ==1'b1) begin 
	o<= 1'b0; 
end

else begin
	if (sel == 1'b0) begin 
		o <= i1;
	end
	else begin
		o <= i2; 
	end 
end 

end

endmodule

`ifdef complex_dsp
module int_sop_2_dspchain (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
	chainin,
	resulta,
	chainout);
input [10:0] mode_sigs;
input clk;
input reset; 
input [17:0] ax, bx;
input [18:0] ay, by;
input [36:0] chainin;

output reg [36:0] resulta;
output reg [36:0] chainout;

int_sop_2 inst1(.clk(clk),.reset(reset),.ax(ax),.bx(bx),.ay(ay),.by(by),.mode_sigs(mode_sigs),.chainin(chainin),.resulta(resulta),.chainout(chainout)); 

endmodule
`else
module int_sop_2_dspchain (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
	chainin,
	resulta,
	chainout);
input [10:0] mode_sigs;
input clk;
input reset; 
input [17:0] ax, bx;
input [18:0] ay, by;
input [36:0] chainin;

output reg [36:0] resulta;
output reg [36:0] chainout;
reg [17:0] ax_reg;
reg [18:0] ay_reg;
reg [17:0] bx_reg;
reg [18:0] by_reg;
reg [36:0] resulta;
always @(posedge clk) begin
  if(reset) begin
    resulta <= 0;
    ax_reg <= 0;
    ay_reg <= 0;
    bx_reg <= 0;
    by_reg <= 0;
  end
  else begin
    ax_reg <= ax;
    ay_reg <= ay;
    bx_reg <= bx;
    by_reg <= by;
    resulta <= ax_reg * ay_reg + bx_reg * by_reg + chainin;
  end
end
assign chainout = resulta;
endmodule
`endif

`ifdef complex_dsp
module fp16_sop2_mult_dspchain (clk,reset,top_a,top_b,bot_a,bot_b,fp32_in,mode_sigs,chainin,chainout,result);
input clk; 
input reset;
input [10:0] mode_sigs; 
input [15:0] top_a,top_b,bot_a,bot_b;
input [31:0] chainin,fp32_in; 
output reg [31:0] chainout, result;

fp16_sop2_mult inst1(.clk(clk),.reset(reset),.top_a(top_a),.top_b(top_b),.bot_a(bot_a),.bot_b(bot_b),.fp32_in(fp32_in),.mode_sigs(mode_sigs),.chainin(chainin),.chainout(chainout),.result(result)); 

endmodule

`else
module fp16_sop2_mult_dspchain (clk,reset,top_a,top_b,bot_a,bot_b,fp32_in,mode_sigs,chainin,chainout,result);
input clk; 
input reset;
input [10:0] mode_sigs; 
input [15:0] top_a,top_b,bot_a,bot_b;
input [31:0] chainin,fp32_in; 
output reg [31:0] chainout, result; 

reg [15:0] top_a_reg,top_b_reg,bot_a_reg,bot_b_reg; 
reg [31:0] chainin_reg; 
reg [31:0] r1,r2,r3; 
always@(posedge clk) begin 
if(reset) begin 
top_a_reg<= 16'b0; 
top_b_reg<= 16'b0; 
bot_a_reg<= 16'b0; 
bot_b_reg<= 16'b0;
//result<=32'b0;
//chainout<=32'b0;
chainin_reg<=32'b0;   
end
else begin 
top_a_reg<=top_a; 
top_b_reg<=top_b; 
bot_a_reg<=bot_a;
bot_b_reg<=bot_b;
//chainout<=result;
chainin_reg<=chainin; 
end
end

wire [4:0] flags1,flags2,flags3,flags4; 

FPMult_16_dspchain inst1(.clk(clk),.rst(reset),.a(top_a_reg),.b(top_b_reg),.flags(flags1),.result(r1)); 
FPMult_16_dspchain inst2(.clk(clk),.rst(reset),.a(bot_a_reg),.b(bot_b_reg),.flags(flags2),.result(r2));
FPAddSub_single_dspchain inst3(.clk(clk),.rst(reset),.a(r1),.b(r2),.flags(flags3),.operation(1'b1),.result(r3));
FPAddSub_single_dspchain inst4(.clk(clk),.rst(reset),.a(r3),.b(chainin),.flags(flags4),.operation(1'b1),.result(result));
assign chainout = result; 
endmodule
//`endif

//`timescale 1ns / 1ps


// IEEE Half Precision => 5 = 5, 10 = 10



//`define IEEE_COMPLIANCE 1


//////////////////////////////////////////////////////////////////////////////////
//
// Module Name:    FPMult
//
//////////////////////////////////////////////////////////////////////////////////

module FPMult_16_dspchain(
		clk,
		rst,
		a,
		b,
		result,
		flags
    );
	
	// Input Ports
	input clk ;							// Clock
	input rst ;							// Reset signal
	input [16-1:0] a;						// Input A, a 32-bit floating point number
	input [16-1:0] b;						// Input B, a 32-bit floating point number
	
	// Output ports
	output [32-1:0] result ;					// Product, result of the operation, 32-bit FP number
	output [4:0] flags ;						// Flags indicating exceptions according to IEEE754
	
	// Internal signals
	wire [32-1:0] Z_int ;					// Product, result of the operation, 32-bit FP number
	wire [4:0] Flags_int ;						// Flags indicating exceptions according to IEEE754
	
	wire Sa ;							// A's sign
	wire Sb ;							// B's sign
	wire Sp ;							// Product sign
	wire [5-1:0] Ea ;					// A's 5
	wire [5-1:0] Eb ;					// B's 5
	wire [2*10+1:0] Mp ;					// Product 10
	wire [4:0] InputExc ;						// Exceptions in inputs
	wire [23-1:0] NormM ;					// Normalized 10
	wire [8:0] NormE ;					// Normalized 5
	wire [23:0] RoundM ;					// Normalized 10
	wire [8:0] RoundE ;					// Normalized 5
	wire [23:0] RoundMP ;					// Normalized 10
	wire [8:0] RoundEP ;					// Normalized 5
	wire GRS ;

	//reg [63:0] pipe_0;						// Pipeline register Input->Prep
	reg [2*16-1:0] pipe_0;					// Pipeline register Input->Prep

	//reg [92:0] pipe_1;						// Pipeline register Prep->Execute
	//reg [3*10+2*5+7:0] pipe_1;			// Pipeline register Prep->Execute
	reg [3*10+2*5+18:0] pipe_1;

	//reg [38:0] pipe_2;						// Pipeline register Execute->Normalize
	reg [23+8+7:0] pipe_2;				// Pipeline register Execute->Normalize

	//reg [72:0] pipe_3;						// Pipeline register Normalize->Round
	reg [2*23+2*8+10:0] pipe_3;			// Pipeline register Normalize->Round

	//reg [36:0] pipe_4;						// Pipeline register Round->Output
	reg [32+4:0] pipe_4;					// Pipeline register Round->Output
	
	assign result = pipe_4[32+4:5] ;
	assign flags = pipe_4[4:0] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPMult_PrepModule_dspchain PrepModule(clk, rst, pipe_0[2*16-1:16], pipe_0[16-1:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10+1:0], InputExc[4:0]) ;

	// Perform (unsigned) 10 multiplication
	FPMult_ExecuteModule_dspchain ExecuteModule(pipe_1[3*10+5*2+7:2*10+2*5+8], pipe_1[2*10+2*5+7:2*10+7], pipe_1[2*10+6:5], pipe_1[2*10+2*5+6:2*10+5+7], pipe_1[2*10+5+6:2*10+7], pipe_1[2*10+2*5+8], pipe_1[2*10+2*5+7], Sp, NormE[8:0], NormM[23-1:0], GRS) ;

	// Round result and if necessary, perform a second (post-rounding) normalization step
	FPMult_NormalizeModule_dspchain NormalizeModule(pipe_2[23-1:0], pipe_2[23+8:23], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]) ;		

	// Round result and if necessary, perform a second (post-rounding) normalization step
	//FPMult_RoundModule RoundModule(pipe_3[47:24], pipe_3[23:0], pipe_3[65:57], pipe_3[56:48], pipe_3[66], pipe_3[67], pipe_3[72:68], Z_int[31:0], Flags_int[4:0]) ;		
	FPMult_RoundModule_dspchain RoundModule(pipe_3[2*23+1:23+1], pipe_3[23:0], pipe_3[2*8+2*23+3:2*23+8+3], pipe_3[2*23+8+2:2*23+2], pipe_3[2*23+2*8+4], pipe_3[2*23+2*8+5], pipe_3[2*23+2*8+10:2*23+2*8+6], Z_int[32-1:0], Flags_int[4:0]) ;		


//adding always@ (*) instead of posedge clock to make design combinational
	always @ (*) begin	
		if(rst) begin
			pipe_0 = 0;
			pipe_1 = 0;
			pipe_2 = 0; 
			pipe_3 = 0;
			pipe_4 = 0;
		end 
		else begin		
			/* PIPE 0
				[2*16-1:16] A
				[16-1:0] B
			*/
                       pipe_0 = {a, b} ;


			/* PIPE 1
				[2*5+3*10 + 18: 2*5+2*10 + 18] //pipe_0[16+10-1:16] , 10 of A
				[2*5+2*10 + 17 :2*5+2*10 + 9] // pipe_0[8:0]
				[2*5+2*10 + 8] Sa
				[2*5+2*10 + 7] Sb
				[2*5+2*10 + 6:5+2*10+7] Ea
				[5 +2*10+6:2*10+7] Eb
				[2*10+1+5:5] Mp
				[4:0] InputExc
			*/
			//pipe_1 <= {pipe_0[16+10-1:16], pipe_0[10_MUL_SPLIT_LSB-1:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10-1:0], InputExc[4:0]} ;
			pipe_1 = {pipe_0[16+10-1:16], pipe_0[8:0], Sa, Sb, Ea[5-1:0], Eb[5-1:0], Mp[2*10+1:0], InputExc[4:0]} ;
			
			/* PIPE 2
				[8 + 23 + 7:8 + 23 + 3] InputExc
				[8 + 23 + 2] GRS
				[8 + 23 + 1] Sp
				[8 + 23:23] NormE
				[23-1:0] NormM
			*/
			pipe_2 = {pipe_1[4:0], GRS, Sp, NormE[8:0], NormM[23-1:0]} ;
			/* PIPE 3
				[2*8+2*23+10:2*8+2*23+6] InputExc
				[2*8+2*23+5] GRS
				[2*8+2*23+4] Sp	
				[2*8+2*23+3:8+2*23+3] RoundE
				[8+2*23+2:2*23+2] RoundEP
				[2*23+1:23+1] RoundM
				[23:0] RoundMP
			*/
			pipe_3 = {pipe_2[8 + 23 + 7:8 + 23 + 1], RoundE[8:0], RoundEP[8:0], RoundM[23:0], RoundMP[23:0]} ;
			/* PIPE 4
				[16+4:5] Z
				[4:0] Flags
			*/				
			pipe_4 = {Z_int[32-1:0], Flags_int[4:0]} ;
		end
	end
		
endmodule



module FPMult_PrepModule_dspchain (
		clk,
		rst,
		a,
		b,
		Sa,
		Sb,
		Ea,
		Eb,
		Mp,
		InputExc
	);
	
	// Input ports
	input clk ;
	input rst ;
	input [16-1:0] a ;								// Input A, a 32-bit floating point number
	input [16-1:0] b ;								// Input B, a 32-bit floating point number
	
	// Output ports
	output Sa ;										// A's sign
	output Sb ;										// B's sign
	output [5-1:0] Ea ;								// A's 5
	output [5-1:0] Eb ;								// B's 5
	output [2*10+1:0] Mp ;							// 10 product
	output [4:0] InputExc ;						// Input numbers are exceptions
	
	// Internal signals							// If signal is high...
	wire ANaN ;										// A is a signalling NaN
	wire BNaN ;										// B is a signalling NaN
	wire AInf ;										// A is infinity
	wire BInf ;										// B is infinity
    wire [10-1:0] Ma;
    wire [10-1:0] Mb;
	
	assign ANaN = &(a[16-2:10]) &  |(a[16-2:10]) ;			// All one 5 and not all zero 10 - NaN
	assign BNaN = &(b[16-2:10]) &  |(b[10-1:0]);			// All one 5 and not all zero 10 - NaN
	assign AInf = &(a[16-2:10]) & ~|(a[16-2:10]) ;		// All one 5 and all zero 10 - Infinity
	assign BInf = &(b[16-2:10]) & ~|(b[16-2:10]) ;		// All one 5 and all zero 10 - Infinity
	
	// Check for any exceptions and put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	//assign InputExc = {(ANaN | ANaN | BNaN |BNaN), ANaN, ANaN, BNaN,BNaN} ;
	
	// Take input numbers apart
	assign Sa = a[16-1] ;							// A's sign
	assign Sb = b[16-1] ;							// B's sign
	assign Ea = a[16-2:10];						// Store A's 5 in Ea, unless A is an exception
	assign Eb = b[16-2:10];						// Store B's 5 in Eb, unless B is an exception	
//    assign Ma = a[10_MSB:10_LSB];
  //  assign Mb = b[10_MSB:10_LSB];
	

	// Actual 10 multiplication occurs here
	//assign Mp = ({4'b0001, a[10-1:0]}*{4'b0001, b[10-1:9]}) ;
	assign Mp = ({1'b1,a[10-1:0]}*{1'b1, b[10-1:0]}) ;

	
    //We multiply part of the 10 here
    //Full 10 of A
    //Bits 10_MUL_SPLIT_MSB:10_MUL_SPLIT_LSB of B
   // wire [`ACTUAL_10-1:0] inp_A;
   // wire [`ACTUAL_10-1:0] inp_B;
   // assign inp_A = {1'b1, Ma};
   // assign inp_B = {{(10-(10_MUL_SPLIT_MSB-10_MUL_SPLIT_LSB+1)){1'b0}}, 1'b1, Mb[10_MUL_SPLIT_MSB:10_MUL_SPLIT_LSB]};
   // DW02_mult #(`ACTUAL_10,`ACTUAL_10) u_mult(.A(inp_A), .B(inp_B), .TC(1'b0), .PRODUCT(Mp));
endmodule


module FPMult_ExecuteModule_dspchain(
		a,
		b,
		MpC,
		Ea,
		Eb,
		Sa,
		Sb,
		Sp,
		NormE,
		NormM,
		GRS
    );

	// Input ports
	input [10-1:0] a ;
	input [2*5:0] b ;
	input [2*10+1:0] MpC ;
	input [5-1:0] Ea ;						// A's 5
	input [5-1:0] Eb ;						// B's 5
	input Sa ;								// A's sign
	input Sb ;								// B's sign
	
	// Output ports
	output Sp ;								// Product sign
	output [8:0] NormE ;													// Normalized 5
	output [23-1:0] NormM ;												// Normalized 10
	output GRS ;
	
	wire [2*10+1:0] Mp ;
	
	assign Sp = (Sa ^ Sb) ;												// Equal signs give a positive product
	
   // wire [`ACTUAL_10-1:0] inp_a;
   // wire [`ACTUAL_10-1:0] inp_b;
   // assign inp_a = {1'b1, a};
   // assign inp_b = {{(10-10_MUL_SPLIT_LSB){1'b0}}, 1'b0, b};
   // DW02_mult #(`ACTUAL_10,`ACTUAL_10) u_mult(.A(inp_a), .B(inp_b), .TC(1'b0), .PRODUCT(Mp_temp));
   // DW01_add #(2*`ACTUAL_10) u_add(.A(Mp_temp), .B(MpC<<10_MUL_SPLIT_LSB), .CI(1'b0), .SUM(Mp), .CO());

	//assign Mp = (MpC<<(2*5+1)) + ({4'b0001, a[10-1:0]}*{1'b0, b[2*5:0]}) ;
	assign Mp = MpC;


	assign NormM = (Mp[2*10+1] ? Mp[2*10:0] : Mp[2*10-1:0]); 	// Check for overflow
	assign NormE = (Ea + Eb + Mp[2*10+1]);								// If so, increment 5
	
	assign GRS = ((Mp[10]&(Mp[10+1]))|(|Mp[10-1:0])) ;
	
endmodule

module FPMult_NormalizeModule_dspchain(
		NormM,
		NormE,
		RoundE,
		RoundEP,
		RoundM,
		RoundMP
    );

	// Input Ports
	input [23-1:0] NormM ;									// Normalized 10
	input [8:0] NormE ;									// Normalized 5

	// Output Ports
	output [8:0] RoundE ;
	output [8:0] RoundEP ;
	output [23:0] RoundM ;
	output [23:0] RoundMP ; 
	
// 5 = 5 
// 5 -1 = 4
// NEED to subtract 2^4 -1 = 15

wire [8-1 : 0] bias;

assign bias =  ((1<< (8 -1)) -1);

	assign RoundE = NormE - 9'd15 - 9'd15 + 9'd127 ;
	assign RoundEP = NormE - 9'd15 - 9'd15 + 9'd127 ;
	assign RoundM = NormM ;
	assign RoundMP = NormM ;

endmodule

module FPMult_RoundModule_dspchain(
		RoundM,
		RoundMP,
		RoundE,
		RoundEP,
		Sp,
		GRS,
		InputExc,
		Z,
		Flags
    );

	// Input Ports
	input [23:0] RoundM ;									// Normalized 10
	input [23:0] RoundMP ;									// Normalized 5
	input [8:0] RoundE ;									// Normalized 10 + 1
	input [8:0] RoundEP ;									// Normalized 5 + 1
	input Sp ;												// Product sign
	input GRS ;
	input [4:0] InputExc ;
	
	// Output Ports
	output [32-1:0] Z ;										// Final product
	output [4:0] Flags ;
	
	// Internal Signals
	wire [8:0] FinalE ;									// Rounded 5
	wire [23:0] FinalM;
	wire [23:0] PreShiftM;
	
	assign PreShiftM = GRS ? RoundMP : RoundM ;	// Round up if R and (G or S)
	
	// Post rounding normalization (potential one bit shift> use shifted 10 if there is overflow)
	assign FinalM = (PreShiftM[23] ? {1'b0, PreShiftM[23:1]} : PreShiftM[23:0]) ;
	assign FinalE = (PreShiftM[23] ? RoundEP : RoundE) ; // Increment 5 if a shift was done
	
	
	assign Z = {Sp, FinalE[8-1:0], FinalM[21-1:0], 2'b0} ;   // Putting the pieces together
	assign Flags = InputExc[4:0];

endmodule


module FPAddSub_single_dspchain(
		clk,
		rst,
		a,
		b,
		operation,
		result,
		flags
	);

// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [31:0] a ;								// Input A, a 32-bit floating point number
	input [31:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [31:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754

	reg [68:0]pipe_1;
	reg [54:0]pipe_2;
	reg [45:0]pipe_3;


//internal module wires

//output ports
	wire Opout;
	wire Sa;
	wire Sb;
	wire MaxAB;
	wire [7:0] CExp;
	wire [4:0] Shift;
	wire [22:0] Mmax;
	wire [4:0] InputExc;
	wire [23:0] Mmin_3;

	wire [32:0] SumS_5 ;
	wire [4:0] Shift_1;							
	wire PSgn ;							
	wire Opr ;	
	
	wire [22:0] NormM ;				// Normalized mantissa
	wire [8:0] NormE ;					// Adjusted exponent
	wire ZeroSum ;						// Zero flag
	wire NegE ;							// Flag indicating negative exponent
	wire R ;								// Round bit
	wire S ;								// Final sticky bit
	wire FG ;

FPAddSub_a_dspchain M1(a,b,operation,Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3);

FpAddSub_b_dspchain M2(pipe_1[51:29],pipe_1[23:0],pipe_1[67],pipe_1[66],pipe_1[65],pipe_1[68],SumS_5,Shift_1,PSgn,Opr);

FPAddSub_c_dspchain M3(pipe_2[54:22],pipe_2[21:17],pipe_2[16:9],NormM,NormE,ZeroSum,NegE,R,S,FG);

FPAddSub_d_dspchain M4(pipe_3[13],pipe_3[22:14],pipe_3[45:23],pipe_3[11],pipe_3[10],pipe_3[9],pipe_3[8],pipe_3[7],pipe_3[6],pipe_3[5],pipe_3[12],pipe_3[4:0],result,flags );


always @ (posedge clk) begin	
		if(rst) begin
			pipe_1 <= 0;
			pipe_2 <= 0;
			pipe_3 <= 0;
		end 
		else begin
/*
pipe_1:
	[68] Opout;
	[67] Sa;
	[66] Sb;
	[65] MaxAB;
	[64:57] CExp;
	[56:52] Shift;
	[51:29] Mmax;
	[28:24] InputExc;
	[23:0] Mmin_3;	
*/

pipe_1 <= {Opout,Sa,Sb,MaxAB,CExp,Shift,Mmax,InputExc,Mmin_3};

/*
pipe_2:
	[54:22]SumS_5;
	[21:17]Shift;
	[16:9]CExp;	
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_2 <= {SumS_5,Shift_1,pipe_1[64:57], pipe_1[67], pipe_1[66], pipe_1[68], pipe_1[65], pipe_1[28:24] };

/*
pipe_3:
	[45:23] NormM ;				
	[22:14] NormE ;					
	[13]ZeroSum ;						
	[12]NegE ;							
	[11]R ;								
	[10]S ;								
	[9]FG ;
	[8]Sa;
	[7]Sb;
	[6]operation;
	[5]MaxAB;	
	[4:0]InputExc
*/

pipe_3 <= {NormM,NormE,ZeroSum,NegE,R,S,FG, pipe_2[8], pipe_2[7], pipe_2[6], pipe_2[5], pipe_2[4:0] };

end
end

endmodule

// Prealign + Align + Shift 1 + Shift 2
module FPAddSub_a_dspchain(
		A,
		B,
		operation,
		Opout,
		Sa,
		Sb,
		MaxAB,
		CExp,
		Shift,
		Mmax,
		InputExc,
		Mmin_3
		
		
	);
	
	// Input ports
	input [31:0] A ;										// Input A, a 32-bit floating point number
	input [31:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	//output ports
	output Opout;
	output Sa;
	output Sb;
	output MaxAB;
	output [7:0] CExp;
	output [4:0] Shift;
	output [22:0] Mmax;
	output [4:0] InputExc;
	output [23:0] Mmin_3;	
							
	wire [9:0] ShiftDet ;							
	wire [30:0] Aout ;
	wire [30:0] Bout ;
	

	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [7:0] DAB ;										// ExpA - ExpB					
	wire [7:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[30:23]) & |(A[22:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[30:23]) & |(B[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[30:23]) & ~|(A[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[30:23]) & ~|(B[22:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
  assign DAB = (A[30:23] + ~(B[30:23]) + 1) ;
	assign DBA = (B[30:23] + ~(A[30:23]) + 1) ;

	assign Sa = A[31] ;									// A's sign bit
	assign Sb = B[31] ;									// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[30:0] ;
	assign Bout = B[30:0] ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Output ports
													// Number of steps to smaller mantissa shift right
	wire [22:0] Mmin_1 ;							// Smaller mantissa 
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (Aout[30:0] < Bout[30:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[9:5] : ShiftDet[4:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin_1 = MaxAB ? Aout[22:0] : Bout[22:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? Bout[22:0]: Aout[22:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? Bout[30:23] : Aout[30:23]) ;	

// Input ports
					// Smaller mantissa after 16|12|8|4 shift
	wire [2:0] Shift_1 ;						// Shift amount
	
	assign Shift_1 = Shift [4:2];

	wire [23:0] Mmin_2 ;						// The smaller mantissa
	
	// Internal signals
	reg	  [23:0]		Lvl1;
	reg	  [23:0]		Lvl2;
	wire    [47:0]    Stage1;	
	integer           i;                // Loop variable
	
	always @(*) begin						
		// Rotate by 16?
		Lvl1 <= Shift_1[2] ? {17'b00000000000000001, Mmin_1[22:16]} : {1'b1, Mmin_1}; 
	end
	
	assign Stage1 = {Lvl1, Lvl1};
	
	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift_1[1:0])
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[23:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[23:19] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[23:15] <= 0; end
			// Rotate by 12	
			2'b11:  begin for (i=0; i<=23; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[23:11] <= 0; end
	  endcase
	end
	
	// Assign output to next shift stage
	assign Mmin_2 = Lvl2;
								// Smaller mantissa after 16|12|8|4 shift
	wire [1:0] Shift_2 ;						// Shift amount
	
	assign Shift_2 =Shift  [1:0] ;
					// The smaller mantissa
	
	// Internal Signal
	reg	  [23:0]		Lvl3;
	wire    [47:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {Mmin_2, Mmin_2};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_2[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[23:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[23] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[23:22] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=23; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[23:21] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin_3 = Lvl3;	

	
endmodule

module FpAddSub_b_dspchain(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		SumS_5,
		Shift,
		PSgn,
		Opr
);
	input [22:0] Mmax ;					// The larger mantissa
	input [23:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	wire [32:0] Sum ;	
						// Output ports
	output [32:0] SumS_5 ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount				// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation

	// Perform effective operation
	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, 8'b00000000} - {Mmin, 8'b00000000}) : ({1'b1, Mmax, 8'b00000000} + {Mmin, 8'b00000000}) ;
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

		// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[32] ? 5'b00000 :	 
		Sum[31] ? 5'b00001 : 
		Sum[30] ? 5'b00010 : 
		Sum[29] ? 5'b00011 : 
		Sum[28] ? 5'b00100 : 
		Sum[27] ? 5'b00101 : 
		Sum[26] ? 5'b00110 : 
		Sum[25] ? 5'b00111 :
		Sum[24] ? 5'b01000 :
		Sum[23] ? 5'b01001 :
		Sum[22] ? 5'b01010 :
		Sum[21] ? 5'b01011 :
		Sum[20] ? 5'b01100 :
		Sum[19] ? 5'b01101 :
		Sum[18] ? 5'b01110 :
		Sum[17] ? 5'b01111 :
		Sum[16] ? 5'b10000 :
		Sum[15] ? 5'b10001 :
		Sum[14] ? 5'b10010 :
		Sum[13] ? 5'b10011 :
		Sum[12] ? 5'b10100 :
		Sum[11] ? 5'b10101 :
		Sum[10] ? 5'b10110 :
		Sum[9] ? 5'b10111 :
		Sum[8] ? 5'b11000 :
		Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [32:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[16:0], 16'b0000000000000000} : Sum; 
	end
	
	// Assign outputs
	assign SumS_5 = Lvl1;	

endmodule

module FPAddSub_c_dspchain(
		SumS_5,
		Shift,
		CExp,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [32:0] SumS_5 ;						// Smaller mantissa after 16|12|8|4 shift
	
	input [4:0] Shift ;						// Shift amount
	
// Input ports
	
	input [7:0] CExp ;
	

	// Output ports
	output [22:0] NormM ;				// Normalized mantissa
	output [8:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;


	wire [3:0]Shift_1;
	assign Shift_1 = Shift [3:0];
	// Output ports
	wire [32:0] SumS_7 ;						// The smaller mantissa
	
	reg	  [32:0]		Lvl2;
	wire    [65:0]    Stage1;	
	reg	  [32:0]		Lvl3;
	wire    [65:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {SumS_5, SumS_5};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[32:0];       		
			// Rotate by 4
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl2[i-33] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift_1[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[32:0];
			// Rotate by 1
			2'b01: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=65; i>=33; i=i-1) begin Lvl3[i-33] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign SumS_7 = Lvl3;						// Take out smaller mantissa



	
	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [8:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [8:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = SumS_7[32] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|SumS_7 ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[8] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = SumS_7[31:9] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = SumS_7[8] ; 
	assign R = SumS_7[7] ;
	assign S = |SumS_7[6:0] ;		
	
endmodule

module FPAddSub_d_dspchain(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		NegE,
		InputExc,
		P,
		Flags 
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [8:0] NormE ;				// Normalized exponent
	input [22:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	

	input NegE ;						// Negative exponent?
	input [4:0] InputExc ;					// Exceptions in inputs A and B

	// Output ports
	output [31:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// 
	wire [31:0] Z ;					// Final result
	wire EOF ;
	
	// Internal signals
	wire [23:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [22:0] RoundM ;				// The final rounded sum
	wire [8:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	wire FSgn;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[22:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[23] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? 8'b00000000 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[7:0], RoundM[22:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[8];

/////////////////////////////////////////////////////////////////////////////////////////////////////////



	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[30:23]) & ~|(Z[30:23]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule

`endif 


module dpram_2048_40bit (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b
);
parameter AWIDTH=11;
parameter NUM_WORDS=2048;
parameter DWIDTH=40;
input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren_a) begin
      ram[address_a] <= data_a;
  end
  else begin
      out_a <= ram[address_a];
  end
end
  
always @ (posedge clk) begin 
  if (wren_b) begin
      ram[address_b] <= data_b;
  end 
  else begin
      out_b <= ram[address_b];
  end
end

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif
endmodule
module dsp_chain_4_fp16_sop2_mult (clk,reset,top_a1,top_b1,bot_a1,bot_b1,top_a2,top_b2,bot_a2,bot_b2,top_a3,top_b3,bot_a3,bot_b3,top_a4,top_b4,bot_a4,bot_b4,result); 

input clk;
input reset; 
input [15:0] top_a1, top_b1, bot_a1, bot_b1, top_a2, top_b2, bot_a2, bot_b2, top_a3, top_b3, bot_a3, bot_b3, top_a4, top_b4, bot_a4, bot_b4; 
output reg [31:0] result; 

wire [31:0] chainin0, chainin1, chainin2, chainin3;
wire [31:0] chainout0, chainout1, chainout2, chainout3; 
wire [31:0] fp32_in1, fp32_in2, fp32_in3, fp32_in4; 
wire [31:0] result1, result2, result3, result4; 

assign fp32_in1 = 32'd0; 
assign fp32_in2 = 32'd0;
assign fp32_in3 = 32'd0;
assign fp32_in4 = 32'd0;
assign chainin0 = 32'd0; 

fp16_sop2_mult_dspchain inst1 (.clk(clk),.reset(reset),.top_a(top_a1),.top_b(top_b1),.bot_a(bot_a1),.bot_b(bot_b1),.fp32_in(fp32_in1),.mode_sigs(11'd0),.chainin(chainin0),.chainout(chainout0),.result(result1)); 
fp16_sop2_mult_dspchain inst2 (.clk(clk),.reset(reset),.top_a(top_a2),.top_b(top_b2),.bot_a(bot_a2),.bot_b(bot_b2),.fp32_in(fp32_in2),.mode_sigs(11'd0),.chainin(chainout0),.chainout(chainout1),.result(result2)); 
fp16_sop2_mult_dspchain inst3 (.clk(clk),.reset(reset),.top_a(top_a3),.top_b(top_b3),.bot_a(bot_a3),.bot_b(bot_b3),.fp32_in(fp32_in3),.mode_sigs(11'd0),.chainin(chainout1),.chainout(chainout2),.result(result3)); 
fp16_sop2_mult_dspchain inst4 (.clk(clk),.reset(reset),.top_a(top_a4),.top_b(top_b4),.bot_a(bot_a4),.bot_b(bot_b4),.fp32_in(fp32_in4),.mode_sigs(11'd0),.chainin(chainout2),.chainout(chainout3),.result(result4)); 

assign result = result4;  


endmodule
module dsp_chain_2_fp16_sop2_mult (clk,reset,top_a1,top_b1,bot_a1,bot_b1,top_a2,top_b2,bot_a2,bot_b2,result); 

input clk;
input reset; 
input [15:0] top_a1, top_b1, bot_a1, bot_b1, top_a2, top_b2, bot_a2, bot_b2; 
output [31:0] result; 

wire [31:0] chainin0, chainin1;
wire [31:0] chainout0, chainout1; 
wire [31:0] fp32_in1, fp32_in2; 
wire [31:0] result1, result2; 

assign fp32_in1 = 32'd0; 
assign fp32_in2 = 32'd0; 
//assign chainin0 = 32'd0; 

fp16_sop2_mult_dspchain inst1 (.clk(clk),.reset(reset),.top_a(top_a1),.top_b(top_b1),.bot_a(bot_a1),.bot_b(bot_b1),.fp32_in(fp32_in1),.mode_sigs(11'd0),.chainin(chainin0),.chainout(chainout0),.result(result1)); 
fp16_sop2_mult_dspchain inst2 (.clk(clk),.reset(reset),.top_a(top_a2),.top_b(top_b2),.bot_a(bot_a2),.bot_b(bot_b2),.fp32_in(fp32_in2),.mode_sigs(11'd0),.chainin(chainout0),.chainout(chainout1),.result(result2)); 

assign result = result2;  


endmodule
module dsp_chain_3_fp16_sop2_mult (clk,reset,top_a1,top_b1,bot_a1,bot_b1,top_a2,top_b2,bot_a2,bot_b2,top_a3,top_b3,bot_a3,bot_b3,result); 

input clk;
input reset; 
input [15:0] top_a1, top_b1, bot_a1, bot_b1, top_a2, top_b2, bot_a2, bot_b2, top_a3, top_b3, bot_a3, bot_b3; 
output reg [31:0] result; 

wire [31:0] chainin0, chainin1, chainin2;
wire [31:0] chainout0, chainout1, chainout2; 
wire [31:0] fp32_in1, fp32_in2, fp32_in3; 
wire [31:0] result1, result2, result3; 

assign fp32_in1 = 32'd0; 
assign fp32_in2 = 32'd0;
assign fp32_in3 = 32'd0;
assign chainin0 = 32'd0; 

fp16_sop2_mult_dspchain inst1 (.clk(clk),.reset(reset),.top_a(top_a1),.top_b(top_b1),.bot_a(bot_a1),.bot_b(bot_b1),.fp32_in(fp32_in1),.mode_sigs(11'd0),.chainin(chainin0),.chainout(chainout0),.result(result1)); 
fp16_sop2_mult_dspchain inst2 (.clk(clk),.reset(reset),.top_a(top_a2),.top_b(top_b2),.bot_a(bot_a2),.bot_b(bot_b2),.fp32_in(fp32_in2),.mode_sigs(11'd0),.chainin(chainout0),.chainout(chainout1),.result(result2)); 
fp16_sop2_mult_dspchain inst3 (.clk(clk),.reset(reset),.top_a(top_a3),.top_b(top_b3),.bot_a(bot_a3),.bot_b(bot_b3),.fp32_in(fp32_in3),.mode_sigs(11'd0),.chainin(chainout1),.chainout(chainout2),.result(result3)); 

assign result = result3;  

endmodule
`define DWIDTH 8
`define DESIGN_SIZE 32
`define MASK_WIDTH 2

module activation_32_8bit(
    input activation_type,
    input enable_activation,
    input in_data_available,
    input [`DESIGN_SIZE*`DWIDTH-1:0] inp_data,
    output [`DESIGN_SIZE*`DWIDTH-1:0] out_data,
    output out_data_available,
    input [`MASK_WIDTH-1:0] validity_mask,
    output done_activation,
    input clk,
    input reset
);

reg  done_activation_internal;
reg  out_data_available_internal;
wire [`DESIGN_SIZE*`DWIDTH-1:0] out_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] slope_applied_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] intercept_applied_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] relu_applied_data_internal;
reg [31:0] i;
reg [31:0] cycle_count;
reg activation_in_progress;

reg [(`DESIGN_SIZE*4)-1:0] address;
reg [(`DESIGN_SIZE*8)-1:0] data_slope;
reg [(`DESIGN_SIZE*8)-1:0] data_slope_flopped;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept_delayed;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept_flopped;

reg in_data_available_flopped;
reg [`DESIGN_SIZE*`DWIDTH-1:0] inp_data_flopped;

always @(posedge clk) begin
  if (reset) begin
    inp_data_flopped <= 0;
    data_slope_flopped <= 0;
  end else begin
    inp_data_flopped <= inp_data;
    data_slope_flopped <= data_slope;
  end
end

// If the activation block is not enabled, just forward the input data
assign out_data             = enable_activation ? out_data_internal : inp_data_flopped;
assign done_activation      = enable_activation ? done_activation_internal : 1'b1;
assign out_data_available   = enable_activation ? out_data_available_internal : in_data_available_flopped;

always @(posedge clk) begin
   if (reset || ~enable_activation) begin
      slope_applied_data_internal     <= 0;
      intercept_applied_data_internal <= 0; 
      relu_applied_data_internal      <= 0; 
      data_intercept_delayed      <= 0;
      data_intercept_flopped      <= 0;
      done_activation_internal    <= 0;
      out_data_available_internal <= 0;
      cycle_count                 <= 0;
      activation_in_progress      <= 0;
      in_data_available_flopped <= in_data_available;
   end else if(in_data_available || activation_in_progress) begin
      cycle_count = cycle_count + 1;

      for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
         if(activation_type==1'b1) begin // tanH
            slope_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= data_slope_flopped[i*8 +: 8] * inp_data_flopped[i*`DWIDTH +:`DWIDTH];
            data_intercept_flopped[i*8 +: 8] <= data_intercept[i*8 +: 8];
            data_intercept_delayed[i*8 +: 8] <= data_intercept_flopped[i*8 +: 8];
            intercept_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= slope_applied_data_internal[i*`DWIDTH +:`DWIDTH] + data_intercept_delayed[i*8 +: 8];
         end else begin // ReLU
            relu_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= inp_data[i*`DWIDTH] ? {`DWIDTH{1'b0}} : inp_data[i*`DWIDTH +:`DWIDTH];
         end
      end   

      //TANH needs 1 extra cycle
      if (activation_type==1'b1) begin
         if (cycle_count==3) begin
            out_data_available_internal <= 1;
         end
      end else begin
         if (cycle_count==2) begin
           out_data_available_internal <= 1;
         end
      end

      //TANH needs 1 extra cycle
      if (activation_type==1'b1) begin
        if(cycle_count==(`DESIGN_SIZE+2)) begin
           done_activation_internal <= 1'b1;
           activation_in_progress <= 0;
        end
        else begin
           activation_in_progress <= 1;
        end
      end else begin
        if(cycle_count==(`DESIGN_SIZE+1)) begin
           done_activation_internal <= 1'b1;
           activation_in_progress <= 0;
        end
        else begin
           activation_in_progress <= 1;
        end
      end
   end
   else begin
      slope_applied_data_internal     <= 0;
      intercept_applied_data_internal <= 0; 
      relu_applied_data_internal      <= 0; 
      data_intercept_delayed      <= 0;
      data_intercept_flopped      <= 0;
      done_activation_internal    <= 0;
      out_data_available_internal <= 0;
      cycle_count                 <= 0;
      activation_in_progress      <= 0;
   end
end

assign out_data_internal = (activation_type) ? intercept_applied_data_internal : relu_applied_data_internal;

//Our equation of tanh is Y=AX+B
//A is the slope and B is the intercept.
//We store A in one LUT and B in another.
//LUT for the slope
always @(address) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
    case (address[i*4+:4])
      4'b0000: data_slope[i*8+:8] = 8'd0;
      4'b0001: data_slope[i*8+:8] = 8'd0;
      4'b0010: data_slope[i*8+:8] = 8'd2;
      4'b0011: data_slope[i*8+:8] = 8'd3;
      4'b0100: data_slope[i*8+:8] = 8'd4;
      4'b0101: data_slope[i*8+:8] = 8'd0;
      4'b0110: data_slope[i*8+:8] = 8'd4;
      4'b0111: data_slope[i*8+:8] = 8'd3;
      4'b1000: data_slope[i*8+:8] = 8'd2;
      4'b1001: data_slope[i*8+:8] = 8'd0;
      4'b1010: data_slope[i*8+:8] = 8'd0;
      default: data_slope[i*8+:8] = 8'd0;
    endcase  
    end
end

//LUT for the intercept
always @(address) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
    case (address[i*4+:4])
      4'b0000: data_intercept[i*8+:8] = 8'd127;
      4'b0001: data_intercept[i*8+:8] = 8'd99;
      4'b0010: data_intercept[i*8+:8] = 8'd46;
      4'b0011: data_intercept[i*8+:8] = 8'd18;
      4'b0100: data_intercept[i*8+:8] = 8'd0;
      4'b0101: data_intercept[i*8+:8] = 8'd0;
      4'b0110: data_intercept[i*8+:8] = 8'd0;
      4'b0111: data_intercept[i*8+:8] = -8'd18;
      4'b1000: data_intercept[i*8+:8] = -8'd46;
      4'b1001: data_intercept[i*8+:8] = -8'd99;
      4'b1010: data_intercept[i*8+:8] = -8'd127;
      default: data_intercept[i*8+:8] = 8'd0;
    endcase  
    end
end

//Logic to find address
always @(inp_data) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
        if((inp_data[i*`DWIDTH +:`DWIDTH])>=90) begin
           address[i*4+:4] = 4'b0000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=39 && (inp_data[i*`DWIDTH +:`DWIDTH])<90) begin
           address[i*4+:4] = 4'b0001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=28 && (inp_data[i*`DWIDTH +:`DWIDTH])<39) begin
           address[i*4+:4] = 4'b0010;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=16 && (inp_data[i*`DWIDTH +:`DWIDTH])<28) begin
           address[i*4+:4] = 4'b0011;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=1 && (inp_data[i*`DWIDTH +:`DWIDTH])<16) begin
           address[i*4+:4] = 4'b0100;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])==0) begin
           address[i*4+:4] = 4'b0101;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-16 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-1) begin
           address[i*4+:4] = 4'b0110;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-28 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-16) begin
           address[i*4+:4] = 4'b0111;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-39 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-28) begin
           address[i*4+:4] = 4'b1000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-90 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-39) begin
           address[i*4+:4] = 4'b1001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])<=-90) begin
           address[i*4+:4] = 4'b1010;
        end
        else begin
           address[i*4+:4] = 4'b0101;
        end
    end
end

//Adding a dummy signal to use validity_mask input, to make ODIN happy
//TODO: Need to correctly use validity_mask
wire [`MASK_WIDTH-1:0] dummy;
assign dummy = validity_mask;

endmodule
`define DWIDTH 16
`define DESIGN_SIZE 32
`define MASK_WIDTH 2

module activation_32_16bit(
    input activation_type,
    input enable_activation,
    input in_data_available,
    input [`DESIGN_SIZE*`DWIDTH-1:0] inp_data,
    output [`DESIGN_SIZE*`DWIDTH-1:0] out_data,
    output out_data_available,
    input [`MASK_WIDTH-1:0] validity_mask,
    output done_activation,
    input clk,
    input reset
);

reg  done_activation_internal;
reg  out_data_available_internal;
wire [`DESIGN_SIZE*`DWIDTH-1:0] out_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] slope_applied_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] intercept_applied_data_internal;
reg [`DESIGN_SIZE*`DWIDTH-1:0] relu_applied_data_internal;
reg [31:0] i;
reg [31:0] cycle_count;
reg activation_in_progress;

reg [(`DESIGN_SIZE*4)-1:0] address;
reg [(`DESIGN_SIZE*8)-1:0] data_slope;
reg [(`DESIGN_SIZE*8)-1:0] data_slope_flopped;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept_delayed;
reg [(`DESIGN_SIZE*8)-1:0] data_intercept_flopped;

reg in_data_available_flopped;
reg [`DESIGN_SIZE*`DWIDTH-1:0] inp_data_flopped;

always @(posedge clk) begin
  if (reset) begin
    inp_data_flopped <= 0;
    data_slope_flopped <= 0;
  end else begin
    inp_data_flopped <= inp_data;
    data_slope_flopped <= data_slope;
  end
end

// If the activation block is not enabled, just forward the input data
assign out_data             = enable_activation ? out_data_internal : inp_data_flopped;
assign done_activation      = enable_activation ? done_activation_internal : 1'b1;
assign out_data_available   = enable_activation ? out_data_available_internal : in_data_available_flopped;

always @(posedge clk) begin
   if (reset || ~enable_activation) begin
      slope_applied_data_internal     <= 0;
      intercept_applied_data_internal <= 0; 
      relu_applied_data_internal      <= 0; 
      data_intercept_delayed      <= 0;
      data_intercept_flopped      <= 0;
      done_activation_internal    <= 0;
      out_data_available_internal <= 0;
      cycle_count                 <= 0;
      activation_in_progress      <= 0;
      in_data_available_flopped <= in_data_available;
   end else if(in_data_available || activation_in_progress) begin
      cycle_count = cycle_count + 1;

      for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
         if(activation_type==1'b1) begin // tanH
            slope_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= data_slope_flopped[i*8 +: 8] * inp_data_flopped[i*`DWIDTH +:`DWIDTH];
            data_intercept_flopped[i*8 +: 8] <= data_intercept[i*8 +: 8];
            data_intercept_delayed[i*8 +: 8] <= data_intercept_flopped[i*8 +: 8];
            intercept_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= slope_applied_data_internal[i*`DWIDTH +:`DWIDTH] + data_intercept_delayed[i*8 +: 8];
         end else begin // ReLU
            relu_applied_data_internal[i*`DWIDTH +:`DWIDTH] <= inp_data[i*`DWIDTH] ? {`DWIDTH{1'b0}} : inp_data[i*`DWIDTH +:`DWIDTH];
         end
      end   

      //TANH needs 1 extra cycle
      if (activation_type==1'b1) begin
         if (cycle_count==3) begin
            out_data_available_internal <= 1;
         end
      end else begin
         if (cycle_count==2) begin
           out_data_available_internal <= 1;
         end
      end

      //TANH needs 1 extra cycle
      if (activation_type==1'b1) begin
        if(cycle_count==(`DESIGN_SIZE+2)) begin
           done_activation_internal <= 1'b1;
           activation_in_progress <= 0;
        end
        else begin
           activation_in_progress <= 1;
        end
      end else begin
        if(cycle_count==(`DESIGN_SIZE+1)) begin
           done_activation_internal <= 1'b1;
           activation_in_progress <= 0;
        end
        else begin
           activation_in_progress <= 1;
        end
      end
   end
   else begin
      slope_applied_data_internal     <= 0;
      intercept_applied_data_internal <= 0; 
      relu_applied_data_internal      <= 0; 
      data_intercept_delayed      <= 0;
      data_intercept_flopped      <= 0;
      done_activation_internal    <= 0;
      out_data_available_internal <= 0;
      cycle_count                 <= 0;
      activation_in_progress      <= 0;
   end
end

assign out_data_internal = (activation_type) ? intercept_applied_data_internal : relu_applied_data_internal;

//Our equation of tanh is Y=AX+B
//A is the slope and B is the intercept.
//We store A in one LUT and B in another.
//LUT for the slope
always @(address) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
    case (address[i*4+:4])
      4'b0000: data_slope[i*8+:8] = 8'd0;
      4'b0001: data_slope[i*8+:8] = 8'd0;
      4'b0010: data_slope[i*8+:8] = 8'd2;
      4'b0011: data_slope[i*8+:8] = 8'd3;
      4'b0100: data_slope[i*8+:8] = 8'd4;
      4'b0101: data_slope[i*8+:8] = 8'd0;
      4'b0110: data_slope[i*8+:8] = 8'd4;
      4'b0111: data_slope[i*8+:8] = 8'd3;
      4'b1000: data_slope[i*8+:8] = 8'd2;
      4'b1001: data_slope[i*8+:8] = 8'd0;
      4'b1010: data_slope[i*8+:8] = 8'd0;
      default: data_slope[i*8+:8] = 8'd0;
    endcase  
    end
end

//LUT for the intercept
always @(address) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
    case (address[i*4+:4])
      4'b0000: data_intercept[i*8+:8] = 8'd127;
      4'b0001: data_intercept[i*8+:8] = 8'd99;
      4'b0010: data_intercept[i*8+:8] = 8'd46;
      4'b0011: data_intercept[i*8+:8] = 8'd18;
      4'b0100: data_intercept[i*8+:8] = 8'd0;
      4'b0101: data_intercept[i*8+:8] = 8'd0;
      4'b0110: data_intercept[i*8+:8] = 8'd0;
      4'b0111: data_intercept[i*8+:8] = -8'd18;
      4'b1000: data_intercept[i*8+:8] = -8'd46;
      4'b1001: data_intercept[i*8+:8] = -8'd99;
      4'b1010: data_intercept[i*8+:8] = -8'd127;
      default: data_intercept[i*8+:8] = 8'd0;
    endcase  
    end
end

//Logic to find address
always @(inp_data) begin
    for (i = 0; i < `DESIGN_SIZE; i=i+1) begin
        if((inp_data[i*`DWIDTH +:`DWIDTH])>=90) begin
           address[i*4+:4] = 4'b0000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=39 && (inp_data[i*`DWIDTH +:`DWIDTH])<90) begin
           address[i*4+:4] = 4'b0001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=28 && (inp_data[i*`DWIDTH +:`DWIDTH])<39) begin
           address[i*4+:4] = 4'b0010;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=16 && (inp_data[i*`DWIDTH +:`DWIDTH])<28) begin
           address[i*4+:4] = 4'b0011;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>=1 && (inp_data[i*`DWIDTH +:`DWIDTH])<16) begin
           address[i*4+:4] = 4'b0100;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])==0) begin
           address[i*4+:4] = 4'b0101;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-16 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-1) begin
           address[i*4+:4] = 4'b0110;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-28 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-16) begin
           address[i*4+:4] = 4'b0111;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-39 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-28) begin
           address[i*4+:4] = 4'b1000;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])>-90 && (inp_data[i*`DWIDTH +:`DWIDTH])<=-39) begin
           address[i*4+:4] = 4'b1001;
        end
        else if ((inp_data[i*`DWIDTH +:`DWIDTH])<=-90) begin
           address[i*4+:4] = 4'b1010;
        end
        else begin
           address[i*4+:4] = 4'b0101;
        end
    end
end

//Adding a dummy signal to use validity_mask input, to make ODIN happy
//TODO: Need to correctly use validity_mask
wire [`MASK_WIDTH-1:0] dummy;
assign dummy = validity_mask;

endmodule
module tanh(
input [15:0] x,
output [15:0] tanh_out);

reg [15:0] lut;
wire [15:0] x_comp;
reg [15:0] tanh_comp;
//reg [15:0] tanh;
reg [4:0] address;


assign x_comp = x[15]? {1'b0,~(x[14:0])}+1'b1:x; // first take 2's complement if x is negative
assign tanh_out = x[15]?(~lut+1'b1):lut; // take 2's complement of tanh if x was negative

always @(address)
begin
  case(address)
  5'd0:  lut =16'b0000100000000010; //address(0.55)
  5'd1:  lut=16'b0000100100100101; //address(0.65)
  5'd2:  lut=16'b0000101000101001; //address(0.75)
  5'd3:  lut=16'b0000101100001110; //address(0.85)
  5'd4:  lut=16'b0000101111010110; //address(0.95)
  5'd5:  lut=16'b0000110010000010; //address(1.05)
  5'd6:  lut=16'b0000110100010101; //address(1.15)
  5'd7:  lut=16'b0000110110010010; //address(1.25)
  5'd8:  lut=16'b0000110111111100; //address(1.35)
  5'd9:  lut=16'b0000111001010100; //address(1.45)
  5'd10:  lut=16'b0000111010011110; //address(1.55)
  5'd11:  lut=16'b0000111011011100; //address(1.65)
  5'd12:  lut=16'b0000111100001111; //address(1.75)
  5'd13:  lut=16'b0000111100111010; //address(1.85)
  5'd14:  lut=16'b0000111101011101; //address(1.95)
  5'd15:  lut=16'b0000111101111010; //address(2.05)
  5'd16:  lut=16'b0000111110010010; //address(2.15)
  5'd17:  lut=16'b0000111110100110; //address(2.25)
  5'd18:  lut=16'b0000111110110110; //address(2.35)
  5'd19:  lut=16'b0000111111000011; //address(2.45)
  5'd20:  lut=16'b0000111111001110; //address(2.55)
  5'd21:  lut=16'b0000111111101011; //address(3.0)
  5'd22:  lut=16'b0001000000000000; //1
  5'd23:  lut=x_comp;
  default: lut=0;
  endcase
end

always@(x)
begin
  /*if(rst == 0)
        tanh_out = 0;
  else
    begin*/
    // first take 2's complement if x is negative
    /*if(x[15] == 1'b1)
        begin
            x_comp = {1'b0,~(x[14:0])}+1'b1;
        end
    else
        begin
            x_comp = x;
    end*/

    // next find the address

    if((x_comp >= 16'h0800) && (x_comp < 16'h3000))
    begin
    case(x_comp[15:12])
        4'b0000:begin
                if((x_comp[11:0] >= 16'h800) && (x_comp[11:0] < 16'h99a))
                    address = 5'd0;
                else if((x_comp[11:0] >= 16'h99a) && (x_comp[11:0] < 16'hb33))
                    address = 5'd1;
                else if((x_comp[11:0] >= 16'hb33) && (x_comp[11:0] < 16'hccd))
                    address = 5'd2;
                else if((x_comp[11:0] >= 16'hccd) && (x_comp[11:0] < 16'he66))
                    address = 5'd3;
                else if(x_comp[11:0] >= 16'he66)
                    address = 5'd4;
                end
        4'b0001:begin
                if((x_comp[11:0] >= 16'h000) && (x_comp[11:0] < 16'h19a))
                    address = 5'd5;
                else if((x_comp[11:0] >= 16'h19a) && (x_comp[11:0] < 16'h333))
                    address = 5'd6;
                else if((x_comp[11:0] >= 16'h333) && (x_comp[11:0] < 16'h4cd))
                    address = 5'd7;
                else if((x_comp[11:0] >= 16'h4cd) && (x_comp[11:0] < 16'h666))
                    address = 5'd8;
                else if((x_comp[11:0] >= 16'h666) && (x_comp[11:0] < 16'h800))
                    address = 5'd9;
                else if((x_comp[11:0] >= 16'h800) && (x_comp[11:0] < 16'h99a))
                    address = 5'd10;
                else if((x_comp[11:0] >= 16'h99a) && (x_comp[11:0] < 16'hb33))
                    address = 5'd11;
                else if((x_comp[11:0] >= 16'hb33) && (x_comp[11:0] < 16'hccd))
                    address = 5'd12;
                else if((x_comp[11:0] >= 16'hccd) && (x_comp[11:0] < 16'he66))
                    address = 5'd13;
                else if(x_comp[11:0] >= 16'he66)
                    address = 5'd14;
                end
        4'b0010:begin
                if((x_comp[11:0] >= 16'h000) && (x_comp[11:0] < 16'h19a))
                    address = 5'd15;
                else if((x_comp[11:0] >= 16'h19a) && (x_comp[11:0] < 16'h333))
                    address = 5'd16;
                else if((x_comp[11:0] >= 16'h333) && (x_comp[11:0] < 16'h4cd))
                    address = 5'd17;
                else if((x_comp[11:0] >= 16'h4cd) && (x_comp[11:0] < 16'h666))
                    address = 5'd18;
                else if((x_comp[11:0] >= 16'h666) && (x_comp[11:0] < 16'h800))
                    address = 5'd19;
                else if((x_comp[11:0] >= 16'h800) && (x_comp[11:0] < 16'h99a))
                    address = 5'd20;
                else if(x_comp[11:0] >= 16'h99a)
                    address = 5'd21;
                end
        default: address = 0;
    endcase
    end

    else if((x_comp >= 16'h0000) && (x_comp < 16'h0800))
           begin
               address = 5'd23;
           end
    else if(x_comp >= 16'h3000)
           begin
               address = 5'd22;
           end
   //end

end


endmodule

module sigmoid(
input [15:0] x,
output [15:0] sig_out
);

reg [15:0] lut;
reg [5:0] address;

assign sig_out = lut;

always @(address)
begin

       case(address)
       6'd0: lut = 16'b0000000000101101; //sig(-4.5)
       6'd1: lut = 16'b0000000000110110; //sig(-4.3)
       6'd2: lut = 16'b0000000001000010; //sig(-4.1)
       6'd3: lut = 16'b0000000001010001; //sig(-3.9)
       6'd4:  lut = 16'b0000000001100010; //sig(-3.7)
       6'd5 :  lut = 16'b0000000001111000; //sig(-3.5)
       6'd6 :  lut= 16'b0000000010010001; //sig(-3.3)
       6'd7 :  lut= 16'b0000000010110000; //sig(-3.1)
       6'd8:  lut= 16'b0000000011010101; //sig(-2.9)
       6'd9 :  lut= 16'b0000000100000010; //sig(-2.7)
       6'd10 :  lut= 16'b0000000100110110; //sig(-2.5)
       6'd11 :  lut= 16'b0000000101110101; //sig(-2.3)
       6'd12 :  lut= 16'b0000000110111110; //sig(-2.1)
       6'd13 :  lut= 16'b0000001000010100; //sig(-1.9)
       6'd14 :  lut= 16'b0000001001111000; //sig(-1.7)
       6'd15 :  lut= 16'b0000001011101011; //sig(-1.5)
       6'd16 :  lut= 16'b0000001101101101; //sig(-1.3)
       6'd17:  lut= 16'b0000001111111110; //sig(-1.1)
       6'd18 :  lut= 16'b0000010010100000; //sig(-0.9)
       6'd19 :  lut= 16'b0000010101001111; //sig(-0.7)
       6'd20 :  lut= 16'b0000011000001010; //sig(-0.5)
       6'd21 :  lut= 16'b0000011011001111; //sig(-0.3)
       6'd22 :  lut= 16'b0000011110011001; //sig(-0.1)
       6'd23 :  lut= 16'b0000100001100110; //sig(0.1)
       6'd24 :  lut= 16'b0000100100110000; //sig(0.3)
       6'd25 :  lut= 16'b0000100111110101; //sig(0.5)
       6'd26 :  lut= 16'b0000101010110000; //sig(0.7)
       6'd27 :  lut= 16'b0000101101100000; //sig(0.9)
       6'd28 :  lut= 16'b0000110000000001; //sig(1.1)
       6'd29 :  lut= 16'b0000110010010010; //sig(1.3)
       6'd30 :  lut= 16'b0000110100010100; //sig(1.5)
       6'd31 :  lut= 16'b0000110110000111; //sig(1.7)
       6'd32 :  lut= 16'b0000110111101011; //sig(1.9)
       6'd33 :  lut= 16'b0000111001000001; //sig(2.1)
       6'd34 :  lut= 16'b0000111010001010; //sig(2.3)
       6'd35 :  lut= 16'b0000111011001001; //sig(2.5)
       6'd36 :  lut= 16'b0000111011111110; //sig(2.7)
       6'd37 :  lut= 16'b0000111100101010; //sig(2.9)
       6'd38 :  lut= 16'b0000111101001111; //sig(3.1)
       6'd39 :  lut= 16'b0000111101101110; //sig(3.3)
       6'd40 :  lut= 16'b0000111110000111; //sig(3.5)
       6'd41 :  lut= 16'b0000111110011101; //sig(3.7)
       6'd42 :  lut= 16'b0000111110101110; //sig(3.9)
       6'd43 :  lut= 16'b0000111110111101; //sig(4.1)
       6'd44 :  lut= 16'b0000111111001001; //sig(4.3)
       6'd45 :  lut= 16'b0000111111010011; //sig(4.5)
       6'd46 :  lut= 16'b0000111111011011; //sig(4.7)
       6'd47 :  lut= 16'b0000000000100100; //sig(-4.7)
       6'd48:   lut= 16'b0000000000000000; //0
       6'd49:   lut= 16'b0001000000000000; //1
       default: lut=0;
        endcase
end


always@(x)
begin

    case({x[15:12]})
        4'b1000:address = 6'd48;
        4'b1001:address = 6'd48;
        4'b1010:address = 6'd48;
        4'b1011:address = 6'd48;
        4'b1100:address = 6'd48;
        4'b1101:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // -3
                    begin
                       address = 6'd8;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address = 6'd9;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address = 6'd10;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd11;
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                        address =  6'd12;
                    end
        4'b1110:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // -2
                    begin
                        address =  6'd13;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address =  6'd14;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address = 6'd15;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd16;
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                        address =  6'd17;
                    end
        4'b1111:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333))  // -1
                    begin
                        address =  6'd18;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address =  6'd19;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address =  6'd20;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd21;                                                                                     
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                        address =  6'd22;
                    end
        4'b0000:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // 0
                    begin
                        address =  6'd23;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address =  6'd24;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address =  6'd25;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd26;
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                        address =  6'd27;
                    end
        4'b0001:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // 1
                    begin
                        address =  6'd28;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                        address =  6'd29;
                    end
                else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                        address =  6'd30;
                    end
                else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                        address =  6'd31;
                    end
                else if(x[11:0] > 12'hccd)
                    begin
                       address =  6'd32;
                    end
        4'b0010:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333))  // 2
                    begin
                      address =  6'd33;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                      address =  6'd34;
                    end
                 else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                       address =  6'd35;
                    end
                 else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                       address =  6'd36;
                    end
                 else if(x[11:0] > 12'hccd)
                    begin
                       address =  6'd37;
                    end
        4'b0011:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) // 3
                    begin
                       address =  6'd38;
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                      address =  6'd39;
                    end
                else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                      address =  6'd40;
                    end
                else if((x[11:0] > 12'h99a) && (x[11:0] <= 12'hccd))
                    begin
                      address = 6'd41;
                    end
               else if(x[11:0] > 12'hccd)
                    begin
                       address = 6'd42;
                    end
        4'b0100:address = 6'd49;
        4'b0101:address = 6'd49;
        4'b0110:address = 6'd49;
        4'b0111:address = 6'd49;
       /* 4'b0100:if((x[11:0] >= 12'h000) && (x[11:0] <= 12'h333)) //4
                    begin
                      address = lut[43];
                    end
                else if((x[11:0] > 12'h333) && (x[11:0] <= 12'h666))
                    begin
                       address = lut[44];
                    end
                else if((x[11:0] > 12'h666) && (x[11:0] <= 12'h99a))
                    begin
                       address = lut[45];
                    end
                else if(x[11:0] > 12'h99a)
                    begin
                        address = lut[46];
                    end
        4'b0101: address = lut[46];
        4'b0110: address = lut[46];
        4'b0111: address = lut[46];  */
        /*default:begin
                        address = 16'h1000;
                end*/
        endcase

end

endmodule

module dpram_4096_40bit (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b
);
parameter AWIDTH=12;
parameter NUM_WORDS=4096;
parameter DWIDTH=40;
input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren_a) begin
      ram[address_a] <= data_a;
  end
  else begin
      out_a <= ram[address_a];
  end
end
  
always @ (posedge clk) begin 
  if (wren_b) begin
      ram[address_b] <= data_b;
  end 
  else begin
      out_b <= ram[address_b];
  end
end

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;


dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif
endmodule
module dpram_4096_60bit (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b
);
parameter AWIDTH=12;
parameter NUM_WORDS=4096;
parameter DWIDTH=60;
input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren_a) begin
      ram[address_a] <= data_a;
  end
  else begin
      out_a <= ram[address_a];
  end
end
  
always @ (posedge clk) begin 
  if (wren_b) begin
      ram[address_b] <= data_b;
  end 
  else begin
      out_b <= ram[address_b];
  end
end

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif
endmodule
module dpram_2048_60bit (
    clk,
    address_a,
    address_b,
    wren_a,
    wren_b,
    data_a,
    data_b,
    out_a,
    out_b
);
parameter AWIDTH=11;
parameter NUM_WORDS=2048;
parameter DWIDTH=60;
input clk;
input [(AWIDTH-1):0] address_a;
input [(AWIDTH-1):0] address_b;
input  wren_a;
input  wren_b;
input [(DWIDTH-1):0] data_a;
input [(DWIDTH-1):0] data_b;
output reg [(DWIDTH-1):0] out_a;
output reg [(DWIDTH-1):0] out_b;

`ifndef hard_mem

reg [DWIDTH-1:0] ram[NUM_WORDS-1:0];
always @ (posedge clk) begin 
  if (wren_a) begin
      ram[address_a] <= data_a;
  end
  else begin
      out_a <= ram[address_a];
  end
end
  
always @ (posedge clk) begin 
  if (wren_b) begin
      ram[address_b] <= data_b;
  end 
  else begin
      out_b <= ram[address_b];
  end
end

`else

defparam u_dual_port_ram.ADDR_WIDTH = AWIDTH;
defparam u_dual_port_ram.DATA_WIDTH = DWIDTH;

dual_port_ram u_dual_port_ram(
.addr1(address_a),
.we1(wren_a),
.data1(data_a),
.out1(out_a),
.addr2(address_b),
.we2(wren_b),
.data2(data_b),
.out2(out_b),
.clk(clk)
);

`endif
endmodule
`define EXPONENT 5
`define MANTISSA 10
`define ACTUAL_MANTISSA 11
`define EXPONENT_LSB 10
`define EXPONENT_MSB 14
`define MANTISSA_LSB 0
`define MANTISSA_MSB 9
`define MANTISSA_MUL_SPLIT_LSB 3
`define MANTISSA_MUL_SPLIT_MSB 9
`define SIGN 1
`define SIGN_LOC 15
`define DWIDTH (`SIGN+`EXPONENT+`MANTISSA)
`define IEEE_COMPLIANCE 1
`define DATAWIDTH 16

module mode4_adder_tree(
  inp0, 
  inp1, 
  inp2, 
  inp3, 
  inp4, 
  inp5, 
  inp6, 
  inp7, 
  mode4_stage0_run,
  mode4_stage1_run,
  mode4_stage2_run,
  mode4_stage3_run,

  clk,
  reset,
  outp
);

  input clk;
  input reset;
  input  [`DATAWIDTH-1 : 0] inp0; 
  input  [`DATAWIDTH-1 : 0] inp1; 
  input  [`DATAWIDTH-1 : 0] inp2; 
  input  [`DATAWIDTH-1 : 0] inp3; 
  input  [`DATAWIDTH-1 : 0] inp4; 
  input  [`DATAWIDTH-1 : 0] inp5; 
  input  [`DATAWIDTH-1 : 0] inp6; 
  input  [`DATAWIDTH-1 : 0] inp7; 
  output [`DATAWIDTH-1 : 0] outp;
  input mode4_stage0_run;
  input mode4_stage1_run;
  input mode4_stage2_run;
  input mode4_stage3_run;

  wire   [`DATAWIDTH-1 : 0] add0_out_stage3;
  reg    [`DATAWIDTH-1 : 0] add0_out_stage3_reg;
  wire   [`DATAWIDTH-1 : 0] add1_out_stage3;
  reg    [`DATAWIDTH-1 : 0] add1_out_stage3_reg;
  wire   [`DATAWIDTH-1 : 0] add2_out_stage3;
  reg    [`DATAWIDTH-1 : 0] add2_out_stage3_reg;
  wire   [`DATAWIDTH-1 : 0] add3_out_stage3;
  reg    [`DATAWIDTH-1 : 0] add3_out_stage3_reg;

  wire   [`DATAWIDTH-1 : 0] add0_out_stage2;
  reg    [`DATAWIDTH-1 : 0] add0_out_stage2_reg;
  wire   [`DATAWIDTH-1 : 0] add1_out_stage2;
  reg    [`DATAWIDTH-1 : 0] add1_out_stage2_reg;

  wire   [`DATAWIDTH-1 : 0] add0_out_stage1;
  reg    [`DATAWIDTH-1 : 0] add0_out_stage1_reg;

  wire   [`DATAWIDTH-1 : 0] add0_out_stage0;
  reg    [`DATAWIDTH-1 : 0] outp;

//  always @(posedge clk) begin
//    if (reset) begin
//      outp <= 0;
//      add0_out_stage3_reg <= 0;
//      add1_out_stage3_reg <= 0;
//      add2_out_stage3_reg <= 0;
//      add3_out_stage3_reg <= 0;
//      add0_out_stage2_reg <= 0;
//      add1_out_stage2_reg <= 0;
//      add0_out_stage1_reg <= 0;
//    end
//
//    if(~reset && mode4_stage3_run) begin
//      add0_out_stage3_reg <= add0_out_stage3;
//      add1_out_stage3_reg <= add1_out_stage3;
//      add2_out_stage3_reg <= add2_out_stage3;
//      add3_out_stage3_reg <= add3_out_stage3;
//    end
//
//    if(~reset && mode4_stage2_run) begin
//      add0_out_stage2_reg <= add0_out_stage2;
//      add1_out_stage2_reg <= add1_out_stage2;
//    end
//
//    if(~reset && mode4_stage1_run) begin
//      add0_out_stage1_reg <= add0_out_stage1;
//    end
//
//    if(~reset && mode4_stage0_run) begin
//      outp <= add0_out_stage0;
//    end
//
//  end


always @ (posedge clk) begin
	if(~reset && mode4_stage3_run) begin
      add0_out_stage3_reg <= add0_out_stage3;
      add1_out_stage3_reg <= add1_out_stage3;
      add2_out_stage3_reg <= add2_out_stage3;
      add3_out_stage3_reg <= add3_out_stage3;
    end
	
	else if (reset) begin
		add0_out_stage3_reg <= 0;
		add1_out_stage3_reg <= 0;
		add2_out_stage3_reg <= 0;
		add3_out_stage3_reg <= 0;
	end
end		

always @ (posedge clk) begin
	if(~reset && mode4_stage2_run) begin
      add0_out_stage2_reg <= add0_out_stage2;
      add1_out_stage2_reg <= add1_out_stage2;
    end
	
	else if (reset) begin
		add0_out_stage2_reg <= 0;
		add1_out_stage2_reg <= 0;
	end
end		

always @ (posedge clk) begin
	if(~reset && mode4_stage1_run) begin
      add0_out_stage1_reg <= add0_out_stage1;
    end
	else if (reset) begin
	add0_out_stage1_reg <= 0;
	end
end

always @ (posedge clk) begin
	if(~reset && mode4_stage0_run) begin
		outp <= add0_out_stage0;
    end
	else if (reset) begin
		outp <= 0;
	end
end	

  wire clk_NC;
  wire rst_NC;
  wire [4:0] flags_NC0, flags_NC1, flags_NC2, flags_NC3;
  wire [4:0] flags_NC4, flags_NC5, flags_NC6, flags_NC7;

  // 0 add, 1 sub
  FPAddSub add0_stage3(.clk(clk), .rst(reset), .a(inp0),	.b(inp1), .operation(1'b0),	.result(add0_out_stage3), .flags(flags_NC0));
  FPAddSub add1_stage3(.clk(clk), .rst(reset), .a(inp2),	.b(inp3), .operation(1'b0),	.result(add1_out_stage3), .flags(flags_NC1));
  FPAddSub add2_stage3(.clk(clk), .rst(reset), .a(inp4),	.b(inp5), .operation(1'b0),	.result(add2_out_stage3), .flags(flags_NC2));
  FPAddSub add3_stage3(.clk(clk), .rst(reset), .a(inp6),	.b(inp7), .operation(1'b0),	.result(add3_out_stage3), .flags(flags_NC3));

  FPAddSub add0_stage2(.clk(clk), .rst(reset), .a(add0_out_stage3_reg),	.b(add1_out_stage3_reg), .operation(1'b0),	.result(add0_out_stage2), .flags(flags_NC4));
  FPAddSub add1_stage2(.clk(clk), .rst(reset), .a(add2_out_stage3_reg),	.b(add3_out_stage3_reg), .operation(1'b0),	.result(add1_out_stage2), .flags(flags_NC5));

  FPAddSub add0_stage1(.clk(clk), .rst(reset), .a(add0_out_stage2_reg),	.b(add1_out_stage2_reg), .operation(1'b0),	.result(add0_out_stage1), .flags(flags_NC6));

  FPAddSub add0_stage0(.clk(clk), .rst(reset), .a(outp),	.b(add0_out_stage1_reg), .operation(1'b0),	.result(add0_out_stage0), .flags(flags_NC7));


//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add0_stage3(.a(inp0),       .b(inp1),      .z(add0_out_stage3), .rnd(3'b000),    .status());
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add1_stage3(.a(inp2),       .b(inp3),      .z(add1_out_stage3), .rnd(3'b000),    .status());
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add2_stage3(.a(inp4),       .b(inp5),      .z(add2_out_stage3), .rnd(3'b000),    .status());
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add3_stage3(.a(inp6),       .b(inp7),      .z(add3_out_stage3), .rnd(3'b000),    .status());
//
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add0_stage2(.a(add0_out_stage3_reg),       .b(add1_out_stage3_reg),      .z(add0_out_stage2), .rnd(3'b000),    .status());
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add1_stage2(.a(add2_out_stage3_reg),       .b(add3_out_stage3_reg),      .z(add1_out_stage2), .rnd(3'b000),    .status());
//
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add0_stage1(.a(add0_out_stage2_reg),       .b(add1_out_stage2_reg),      .z(add0_out_stage1), .rnd(3'b000),    .status());
//
//  DW_fp_add #(`MANTISSA, `EXPONENT, `IEEE_COMPLIANCE) add0_stage0(.a(outp),       .b(add0_out_stage1_reg),      .z(add0_out_stage0), .rnd(3'b000),    .status());

endmodule

module FPAddSub(
		clk,
		rst,
		a,
		b,
		operation,			// 0 add, 1 sub
		result,
		flags
	);
	
	// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [`DWIDTH-1:0] a ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [`DWIDTH-1:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754
	
	assign flags = 5'b0;
	
//`ifdef complex_dsp
//adder_fp_clk u_add(.clk(clk), .a(a), .b(b),.out(result));
//`else
FPAddSub_16 u_FPAddSub (.clk(clk), .rst(rst), .a(a), .b(b), .operation(1'b0), .result(result), .flags());
//`endif
endmodule

module FPAddSub_16(
		//bf16,
		clk,
		rst,
		a,
		b,
		operation,			// 0 add, 1 sub
		result,
		flags
	);
	//input bf16; //1 for Bfloat16, 0 for IEEE half precision

	// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [`DWIDTH-1:0] a ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [`DWIDTH-1:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754
	
	// Pipeline Registers
	//reg [79:0] pipe_1;							// Pipeline register PreAlign->Align1
	reg [2*`EXPONENT + 2*`DWIDTH + 5:0] pipe_1;							// Pipeline register PreAlign->Align1

	//reg [67:0] pipe_2;							// Pipeline register Align1->Align3
	//reg [2*`EXPONENT+ 2*`MANTISSA + 8:0] pipe_2;							// Pipeline register Align1->Align3
	wire [2*`EXPONENT+ 2*`MANTISSA + 8:0] pipe_2;

	//reg [76:0] pipe_3;	68						// Pipeline register Align1->Align3
	reg [2*`EXPONENT+ 2*`MANTISSA + 9:0] pipe_3;							// Pipeline register Align1->Align3

	//reg [69:0] pipe_4;							// Pipeline register Align3->Execute
	//reg [2*`EXPONENT+ 2*`MANTISSA + 9:0] pipe_4;							// Pipeline register Align3->Execute
	wire [2*`EXPONENT+ 2*`MANTISSA + 9:0] pipe_4;
	
	//reg [51:0] pipe_5;							// Pipeline register Execute->Normalize
	reg [`DWIDTH+`EXPONENT+11:0] pipe_5;							// Pipeline register Execute->Normalize

	//reg [56:0] pipe_6;							// Pipeline register Nomalize->NormalizeShift1
	//reg [`DWIDTH+`EXPONENT+16:0] pipe_6;							// Pipeline register Nomalize->NormalizeShift1
	wire [`DWIDTH+`EXPONENT+16:0] pipe_6;

	//reg [56:0] pipe_7;							// Pipeline register NormalizeShift2->NormalizeShift3
	//reg [`DWIDTH+`EXPONENT+16:0] pipe_7;							// Pipeline register NormalizeShift2->NormalizeShift3
	wire [`DWIDTH+`EXPONENT+16:0] pipe_7;
	//reg [54:0] pipe_8;							// Pipeline register NormalizeShift3->Round
	reg [`EXPONENT*2+`MANTISSA+15:0] pipe_8;							// Pipeline register NormalizeShift3->Round

	//reg [40:0] pipe_9;							// Pipeline register NormalizeShift3->Round
	//reg [`DWIDTH+8:0] pipe_9;							// Pipeline register NormalizeShift3->Round
	wire [`DWIDTH+8:0] pipe_9;

	// Internal wires between modules
	wire [`DWIDTH-2:0] Aout_0 ;							// A - sign
	wire [`DWIDTH-2:0] Bout_0 ;							// B - sign
	wire Opout_0 ;									// A's sign
	wire Sa_0 ;										// A's sign
	wire Sb_0 ;										// B's sign
	wire MaxAB_1 ;									// Indicates the larger of A and B(0/A, 1/B)
	wire [`EXPONENT-1:0] CExp_1 ;							// Common Exponent
	wire [`EXPONENT-1:0] Shift_1 ;							// Number of steps to smaller mantissa shift right (align)
	wire [`MANTISSA-1:0] Mmax_1 ;							// Larger mantissa
	wire [4:0] InputExc_0 ;						// Input numbers are exceptions
	wire [2*`EXPONENT-1:0] ShiftDet_0 ;
	wire [`MANTISSA-1:0] MminS_1 ;						// Smaller mantissa after 0/16 shift
	wire [`MANTISSA:0] MminS_2 ;						// Smaller mantissa after 0/4/8/12 shift
	wire [`MANTISSA:0] Mmin_3 ;							// Smaller mantissa after 0/1/2/3 shift
	wire [`DWIDTH:0] Sum_4 ;
	wire PSgn_4 ;
	wire Opr_4 ;
	wire [`EXPONENT-1:0] Shift_5 ;							// Number of steps to shift sum left (normalize)
	wire [`DWIDTH:0] SumS_5 ;							// Sum after 0/16 shift
	wire [`DWIDTH:0] SumS_6 ;							// Sum after 0/16 shift
	wire [`DWIDTH:0] SumS_7 ;							// Sum after 0/16 shift
	wire [`MANTISSA-1:0] NormM_8 ;						// Normalized mantissa
	wire [`EXPONENT:0] NormE_8;							// Adjusted exponent
	wire ZeroSum_8 ;								// Zero flag
	wire NegE_8 ;									// Flag indicating negative exponent
	wire R_8 ;										// Round bit
	wire S_8 ;										// Final sticky bit
	wire FG_8 ;										// Final sticky bit
	wire [`DWIDTH-1:0] P_int ;
	wire EOF ;
	
	// Prepare the operands for alignment and check for exceptions
	FPAddSub_PrealignModule PrealignModule
	(	// Inputs
		a, b, operation,
		// Outputs
		Sa_0, Sb_0, ShiftDet_0[2*`EXPONENT-1:0], InputExc_0[4:0], Aout_0[`DWIDTH-2:0], Bout_0[`DWIDTH-2:0], Opout_0) ;
		
	// Prepare the operands for alignment and check for exceptions
	FPAddSub_AlignModule AlignModule
	(	// Inputs
		pipe_1[2*`EXPONENT + 2*`DWIDTH + 4: 2*`EXPONENT +`DWIDTH + 6], pipe_1[2*`EXPONENT +`DWIDTH + 5 :  2*`EXPONENT +7], pipe_1[2*`EXPONENT+4:5],
		// Outputs
		CExp_1[`EXPONENT-1:0], MaxAB_1, Shift_1[`EXPONENT-1:0], MminS_1[`MANTISSA-1:0], Mmax_1[`MANTISSA-1:0]) ;	

	// Alignment Shift Stage 1
	FPAddSub_AlignShift1 AlignShift1
	(  // Inputs
		//bf16, 
		pipe_2[`MANTISSA-1:0], pipe_2[`EXPONENT+ 2*`MANTISSA + 4 : 2*`MANTISSA + 7],
		// Outputs
		MminS_2[`MANTISSA:0]) ;

	// Alignment Shift Stage 3 and compution of guard and sticky bits
	FPAddSub_AlignShift2 AlignShift2  
	(  // Inputs
		pipe_3[`MANTISSA:0], pipe_3[2*`MANTISSA+7:2*`MANTISSA+6],
		// Outputs
		Mmin_3[`MANTISSA:0]) ;
						
	// Perform mantissa addition
	FPAddSub_ExecutionModule ExecutionModule
	(  // Inputs
		pipe_4[`MANTISSA*2+5:`MANTISSA+6], pipe_4[`MANTISSA:0], pipe_4[2*`EXPONENT+ 2*`MANTISSA + 8], pipe_4[2*`EXPONENT+ 2*`MANTISSA + 7], pipe_4[2*`EXPONENT+ 2*`MANTISSA + 6], pipe_4[2*`EXPONENT+ 2*`MANTISSA + 9],
		// Outputs
		Sum_4[`DWIDTH:0], PSgn_4, Opr_4) ;
	
	// Prepare normalization of result
	FPAddSub_NormalizeModule NormalizeModule
	(  // Inputs
		pipe_5[`DWIDTH:0], 
		// Outputs
		SumS_5[`DWIDTH:0], Shift_5[4:0]) ;
					
	// Normalization Shift Stage 1
	FPAddSub_NormalizeShift1 NormalizeShift1
	(  // Inputs
		pipe_6[`DWIDTH:0], pipe_6[`DWIDTH+`EXPONENT+14:`DWIDTH+`EXPONENT+11],
		// Outputs
		SumS_7[`DWIDTH:0]) ;
		
	// Normalization Shift Stage 3 and final guard, sticky and round bits
	FPAddSub_NormalizeShift2 NormalizeShift2
	(  // Inputs
		pipe_7[`DWIDTH:0], pipe_7[`DWIDTH+`EXPONENT+5:`DWIDTH+6], pipe_7[`DWIDTH+`EXPONENT+15:`DWIDTH+`EXPONENT+11],
		// Outputs
		NormM_8[`MANTISSA-1:0], NormE_8[`EXPONENT:0], ZeroSum_8, NegE_8, R_8, S_8, FG_8) ;

	// Round and put result together
	FPAddSub_RoundModule RoundModule
	(  // Inputs
		 pipe_8[3], pipe_8[4+`EXPONENT:4], pipe_8[`EXPONENT+`MANTISSA+4:5+`EXPONENT], pipe_8[1], pipe_8[0], pipe_8[`EXPONENT*2+`MANTISSA+15], pipe_8[`EXPONENT*2+`MANTISSA+12], pipe_8[`EXPONENT*2+`MANTISSA+11], pipe_8[`EXPONENT*2+`MANTISSA+14], pipe_8[`EXPONENT*2+`MANTISSA+10], 
		// Outputs
		P_int[`DWIDTH-1:0], EOF) ;
	
	// Check for exceptions
	FPAddSub_ExceptionModule Exceptionmodule
	(  // Inputs
		pipe_9[8+`DWIDTH:9], pipe_9[8], pipe_9[7], pipe_9[6], pipe_9[5:1], pipe_9[0], 
		// Outputs
		result[`DWIDTH-1:0], flags[4:0]) ;			
	

assign pipe_2 = {pipe_1[2*`EXPONENT + 2*`DWIDTH + 5], pipe_1[2*`EXPONENT +6:2*`EXPONENT +5], MaxAB_1, CExp_1[`EXPONENT-1:0], Shift_1[`EXPONENT-1:0], Mmax_1[`MANTISSA-1:0], pipe_1[4:0], MminS_1[`MANTISSA-1:0]} ;
assign pipe_4 = {pipe_3[2*`EXPONENT+ 2*`MANTISSA + 9:`MANTISSA+1], Mmin_3[`MANTISSA:0]} ;
assign pipe_6 = {pipe_5[`DWIDTH+`EXPONENT+11], Shift_5[4:0], pipe_5[`DWIDTH+`EXPONENT+10:`DWIDTH+1], SumS_5[`DWIDTH:0]} ;
assign pipe_7 = {pipe_6[`DWIDTH+`EXPONENT+16:`DWIDTH+1], SumS_7[`DWIDTH:0]} ;
assign pipe_9 = {P_int[`DWIDTH-1:0], pipe_8[2], pipe_8[1], pipe_8[0], pipe_8[`EXPONENT+`MANTISSA+9:`EXPONENT+`MANTISSA+5], EOF} ;

	always @ (posedge clk) begin	
		if(rst) begin
			pipe_1 <= 0;
			//pipe_2 <= 0;
			pipe_3 <= 0;
			//pipe_4 <= 0;
			pipe_5 <= 0;
			//pipe_6 <= 0;
			//pipe_7 <= 0;
			pipe_8 <= 0;
			//pipe_9 <= 0;
		end 
		else begin
/* PIPE_1:
	[2*`EXPONENT + 2*`DWIDTH + 5]  Opout_0
	[2*`EXPONENT + 2*`DWIDTH + 4: 2*`EXPONENT +`DWIDTH + 6] A_out0
	[2*`EXPONENT +`DWIDTH + 5 :  2*`EXPONENT +7] Bout_0
	[2*`EXPONENT +6] Sa_0
	[2*`EXPONENT +5] Sb_0
	[2*`EXPONENT +4 : 5] ShiftDet_0
	[4:0] Input Exc
*/
			pipe_1 <= {Opout_0, Aout_0[`DWIDTH-2:0], Bout_0[`DWIDTH-2:0], Sa_0, Sb_0, ShiftDet_0[2*`EXPONENT -1:0], InputExc_0[4:0]} ;	
/* PIPE_2
[2*`EXPONENT+ 2*`MANTISSA + 8] operation
[2*`EXPONENT+ 2*`MANTISSA + 7] Sa_0
[2*`EXPONENT+ 2*`MANTISSA + 6] Sb_0
[2*`EXPONENT+ 2*`MANTISSA + 5] MaxAB_0
[2*`EXPONENT+ 2*`MANTISSA + 4:`EXPONENT+ 2*`MANTISSA + 5] CExp_0
[`EXPONENT+ 2*`MANTISSA + 4 : 2*`MANTISSA + 5] Shift_0
[2*`MANTISSA + 4:`MANTISSA + 5] Mmax_0
[`MANTISSA + 4 : `MANTISSA] InputExc_0
[`MANTISSA-1:0] MminS_1
*/
			//pipe_2 <= {pipe_1[2*`EXPONENT + 2*`DWIDTH + 5], pipe_1[2*`EXPONENT +6:2*`EXPONENT +5], MaxAB_1, CExp_1[`EXPONENT-1:0], Shift_1[`EXPONENT-1:0], Mmax_1[`MANTISSA-1:0], pipe_1[4:0], MminS_1[`MANTISSA-1:0]} ;	
/* PIPE_3
[2*`EXPONENT+ 2*`MANTISSA + 9] operation
[2*`EXPONENT+ 2*`MANTISSA + 8] Sa_0
[2*`EXPONENT+ 2*`MANTISSA + 7] Sb_0
[2*`EXPONENT+ 2*`MANTISSA + 6] MaxAB_0
[2*`EXPONENT+ 2*`MANTISSA + 5:`EXPONENT+ 2*`MANTISSA + 6] CExp_0
[`EXPONENT+ 2*`MANTISSA + 5 : 2*`MANTISSA + 6] Shift_0
[2*`MANTISSA + 5:`MANTISSA + 6] Mmax_0
[`MANTISSA + 5 : `MANTISSA + 1] InputExc_0
[`MANTISSA:0] MminS_2
*/
			pipe_3 <= {pipe_2[2*`EXPONENT+ 2*`MANTISSA + 8:`MANTISSA], MminS_2[`MANTISSA:0]} ;	
/* PIPE_4
[2*`EXPONENT+ 2*`MANTISSA + 9] operation
[2*`EXPONENT+ 2*`MANTISSA + 8] Sa_0
[2*`EXPONENT+ 2*`MANTISSA + 7] Sb_0
[2*`EXPONENT+ 2*`MANTISSA + 6] MaxAB_0
[2*`EXPONENT+ 2*`MANTISSA + 5:`EXPONENT+ 2*`MANTISSA + 6] CExp_0
[`EXPONENT+ 2*`MANTISSA + 5 : 2*`MANTISSA + 6] Shift_0
[2*`MANTISSA + 5:`MANTISSA + 6] Mmax_0
[`MANTISSA + 5 : `MANTISSA + 1] InputExc_0
[`MANTISSA:0] MminS_3
*/				
			//pipe_4 <= {pipe_3[2*`EXPONENT+ 2*`MANTISSA + 9:`MANTISSA+1], Mmin_3[`MANTISSA:0]} ;	
/* PIPE_5 :
[`DWIDTH+ `EXPONENT + 11] operation
[`DWIDTH+ `EXPONENT + 10] PSgn_4
[`DWIDTH+ `EXPONENT + 9] Opr_4
[`DWIDTH+ `EXPONENT + 8] Sa_0
[`DWIDTH+ `EXPONENT + 7] Sb_0
[`DWIDTH+ `EXPONENT + 6] MaxAB_0
[`DWIDTH+ `EXPONENT + 5 :`DWIDTH+6] CExp_0
[`DWIDTH+5:`DWIDTH+1] InputExc_0
[`DWIDTH:0] Sum_4
*/					
			pipe_5 <= {pipe_4[2*`EXPONENT+ 2*`MANTISSA + 9], PSgn_4, Opr_4, pipe_4[2*`EXPONENT+ 2*`MANTISSA + 8:`EXPONENT+ 2*`MANTISSA + 6], pipe_4[`MANTISSA+5:`MANTISSA+1], Sum_4[`DWIDTH:0]} ;
/* PIPE_6 :
[`DWIDTH+ `EXPONENT + 16] operation
[`DWIDTH+ `EXPONENT + 15:`DWIDTH+ `EXPONENT + 11] Shift_5
[`DWIDTH+ `EXPONENT + 10] PSgn_4
[`DWIDTH+ `EXPONENT + 9] Opr_4
[`DWIDTH+ `EXPONENT + 8] Sa_0
[`DWIDTH+ `EXPONENT + 7] Sb_0
[`DWIDTH+ `EXPONENT + 6] MaxAB_0
[`DWIDTH+ `EXPONENT + 5 :`DWIDTH+6] CExp_0
[`DWIDTH+5:`DWIDTH+1] InputExc_0
[`DWIDTH:0] Sum_4
*/				
			//pipe_6 <= {pipe_5[`DWIDTH+`EXPONENT+11], Shift_5[4:0], pipe_5[`DWIDTH+`EXPONENT+10:`DWIDTH+1], SumS_5[`DWIDTH:0]} ;	
/* PIPE_7 :
[`DWIDTH+ `EXPONENT + 16] operation
[`DWIDTH+ `EXPONENT + 15:`DWIDTH+ `EXPONENT + 11] Shift_5
[`DWIDTH+ `EXPONENT + 10] PSgn_4
[`DWIDTH+ `EXPONENT + 9] Opr_4
[`DWIDTH+ `EXPONENT + 8] Sa_0
[`DWIDTH+ `EXPONENT + 7] Sb_0
[`DWIDTH+ `EXPONENT + 6] MaxAB_0
[`DWIDTH+ `EXPONENT + 5 :`DWIDTH+6] CExp_0
[`DWIDTH+5:`DWIDTH+1] InputExc_0
[`DWIDTH:0] Sum_4
*/						
			//pipe_7 <= {pipe_6[`DWIDTH+`EXPONENT+16:`DWIDTH+1], SumS_7[`DWIDTH:0]} ;	
/* PIPE_8:
[2*`EXPONENT + `MANTISSA + 15] FG_8 
[2*`EXPONENT + `MANTISSA + 14] operation
[2*`EXPONENT + `MANTISSA + 13] PSgn_4
[2*`EXPONENT + `MANTISSA + 12] Sa_0
[2*`EXPONENT + `MANTISSA + 11] Sb_0
[2*`EXPONENT + `MANTISSA + 10] MaxAB_0
[2*`EXPONENT + `MANTISSA + 9:`EXPONENT + `MANTISSA + 10] CExp_0
[`EXPONENT + `MANTISSA + 9:`EXPONENT + `MANTISSA + 5] InputExc_8
[`EXPONENT + `MANTISSA + 4 :`EXPONENT + 5] NormM_8 
[`EXPONENT + 4 :4] NormE_8
[3] ZeroSum_8
[2] NegE_8
[1] R_8
[0] S_8
*/				
			pipe_8 <= {FG_8, pipe_7[`DWIDTH+`EXPONENT+16], pipe_7[`DWIDTH+`EXPONENT+10], pipe_7[`DWIDTH+`EXPONENT+8:`DWIDTH+1], NormM_8[`MANTISSA-1:0], NormE_8[`EXPONENT:0], ZeroSum_8, NegE_8, R_8, S_8} ;	
/* pipe_9:
[`DWIDTH + 8 :9] P_int
[8] NegE_8
[7] R_8
[6] S_8
[5:1] InputExc_8
[0] EOF
*/				
			//pipe_9 <= {P_int[`DWIDTH-1:0], pipe_8[2], pipe_8[1], pipe_8[0], pipe_8[`EXPONENT+`MANTISSA+9:`EXPONENT+`MANTISSA+5], EOF} ;	
		end
	end		
	
endmodule


//
// Description:	 	The pre-alignment module is responsible for taking the inputs
//							apart and checking the parts for exceptions.
//							The exponent difference is also calculated in this module.
//


module FPAddSub_PrealignModule(
		A,
		B,
		operation,
		Sa,
		Sb,
		ShiftDet,
		InputExc,
		Aout,
		Bout,
		Opout
	);
	
	// Input ports
	input [`DWIDTH-1:0] A ;										// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	// Output ports
	output Sa ;												// A's sign
	output Sb ;												// B's sign
	output [2*`EXPONENT-1:0] ShiftDet ;
	output [4:0] InputExc ;								// Input numbers are exceptions
	output [`DWIDTH-2:0] Aout ;
	output [`DWIDTH-2:0] Bout ;
	output Opout ;
	
	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [`EXPONENT-1:0] DAB ;										// ExpA - ExpB					
	wire [`EXPONENT-1:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & |(A[`MANTISSA-1:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & |(B[`MANTISSA-1:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & ~|(A[`MANTISSA-1:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & ~|(B[`MANTISSA-1:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
	assign DAB = (A[`DWIDTH-2:`MANTISSA] + ~(B[`DWIDTH-2:`MANTISSA]) + 1) ;
	assign DBA = (B[`DWIDTH-2:`MANTISSA] + ~(A[`DWIDTH-2:`MANTISSA]) + 1) ;
	
	assign Sa = A[`DWIDTH-1] ;									// A's sign bit
	assign Sb = B[`DWIDTH-1] ;									// B's sign	bit
	assign ShiftDet = {DBA[`EXPONENT-1:0], DAB[`EXPONENT-1:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[`DWIDTH-2:0] ;
	assign Bout = B[`DWIDTH-2:0] ;
	
endmodule


//
// Description:	 	The alignment module determines the larger input operand and
//							sets the mantissas, shift and common exponent accordingly.
//


module FPAddSub_AlignModule (
		A,
		B,
		ShiftDet,
		CExp,
		MaxAB,
		Shift,
		Mmin,
		Mmax
	);
	
	// Input ports
	input [`DWIDTH-2:0] A ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-2:0] B ;								// Input B, a 32-bit floating point number
	input [2*`EXPONENT-1:0] ShiftDet ;
	
	// Output ports
	output [`EXPONENT-1:0] CExp ;							// Common Exponent
	output MaxAB ;									// Incidates larger of A and B (0/A, 1/B)
	output [`EXPONENT-1:0] Shift ;							// Number of steps to smaller mantissa shift right
	output [`MANTISSA-1:0] Mmin ;							// Smaller mantissa 
	output [`MANTISSA-1:0] Mmax ;							// Larger mantissa
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (A[`DWIDTH-2:0] < B[`DWIDTH-2:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[2*`EXPONENT-1:`EXPONENT] : ShiftDet[`EXPONENT-1:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin = MaxAB ? A[`MANTISSA-1:0] : B[`MANTISSA-1:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? B[`MANTISSA-1:0]: A[`MANTISSA-1:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? B[`MANTISSA+`EXPONENT-1:`MANTISSA] : A[`MANTISSA+`EXPONENT-1:`MANTISSA]) ;		
	
endmodule


// Description:	 Alignment shift stage 1, performs 16|12|8|4 shift
//


// ONLY THIS MODULE IS HARDCODED for half precision fp16 and bfloat16
module FPAddSub_AlignShift1(
		//bf16,
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	//input bf16;
	input [`MANTISSA-1:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [`EXPONENT-3:0] Shift ;						// Shift amount. Last 2 bits of shifting are done in next stage. Hence, we have [`EXPONENT - 2] bits
	
	// Output ports
	output [`MANTISSA:0] Mmin ;						// The smaller mantissa
	

	wire bf16;
	assign bf16 = 1'b1; //hardcoding to 1, to avoid ODIN issue. a `ifdef here wasn't working. apparently, nested `ifdefs don't work

	// Internal signals
	reg	  [`MANTISSA:0]		Lvl1;
	reg	  [`MANTISSA:0]		Lvl2;
	wire    [2*`MANTISSA+1:0]    Stage1;	
	integer           i;                // Loop variable

	wire [`MANTISSA:0] temp_0; 

assign temp_0 = 0;

	always @(*) begin
		if (bf16 == 1'b1) begin						
//hardcoding for bfloat16
	//For bfloat16, we can shift the mantissa by a max of 7 bits since mantissa has a width of 7. 
	//Hence if either, bit[3]/bit[4]/bit[5]/bit[6]/bit[7] is 1, we can make it 0. This corresponds to bits [5:1] in our updated shift which doesn't contain last 2 bits.
		//Lvl1 <= (Shift[1]|Shift[2]|Shift[3]|Shift[4]|Shift[5]) ? {temp_0} : {1'b1, MminP};  // MANTISSA + 1 width	
		Lvl1 <= (|Shift[`EXPONENT-3:1]) ? {temp_0} : {1'b1, MminP};  // MANTISSA + 1 width	
		end
		else begin
		//for half precision fp16, 10 bits can be shifted. Hence, only shifts till 10 (01010)can be made. 
		Lvl1 <= Shift[2] ? {temp_0} : {1'b1, MminP};
		end
	end
	
	assign Stage1 = { temp_0, Lvl1}; //2*MANTISSA + 2 width

	always @(*) begin    					// Rotate {0 | 4 } bits
	if(bf16 == 1'b1) begin
	  case (Shift[0])
			// Rotate by 0	
			1'b0:  Lvl2 <= Stage1[`MANTISSA:0];       			
			// Rotate by 4	
			1'b1:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[`MANTISSA:`MANTISSA-3] <= 0; end
	  endcase
	end
	else begin
	  case (Shift[1:0])					// Rotate {0 | 4 | 8} bits
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[`MANTISSA:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end Lvl2[`MANTISSA:`MANTISSA-3] <= 0; end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end Lvl2[`MANTISSA:`MANTISSA-7] <= 0; end
			// Rotate by 12	
			2'b11: Lvl2[`MANTISSA: 0] <= 0; 
			//2'b11:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[`MANTISSA:`MANTISSA-12] <= 0; end
	  endcase
	end
	end

	// Assign output to next shift stage
	assign Mmin = Lvl2;
	
endmodule


// Description:	 Alignment shift stage 2, performs 3|2|1 shift
//


module FPAddSub_AlignShift2(
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	input [`MANTISSA:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [1:0] Shift ;						// Shift amount. Last 2 bits
	
	// Output ports
	output [`MANTISSA:0] Mmin ;						// The smaller mantissa
	
	// Internal Signal
	reg	  [`MANTISSA:0]		Lvl3;
	wire    [2*`MANTISSA+1:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {11'b0, MminP};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[`MANTISSA:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end Lvl3[`MANTISSA] <= 0; end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end Lvl3[`MANTISSA:`MANTISSA-1] <= 0; end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end Lvl3[`MANTISSA:`MANTISSA-2] <= 0; end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin = Lvl3;						// Take out smaller mantissa				

endmodule


//
// Description:	 Module that executes the addition or subtraction on mantissas.
//


module FPAddSub_ExecutionModule(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		Sum,
		PSgn,
		Opr
    );

	// Input ports
	input [`MANTISSA-1:0] Mmax ;					// The larger mantissa
	input [`MANTISSA:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	output [`DWIDTH:0] Sum ;					// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	wire [`EXPONENT-1:0]temp_1;

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation
	assign temp_1 = 0;
	// Perform effective operation
//SAMIDH_UNSURE 5--> 8

	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, temp_1} - {Mmin, temp_1}) : ({1'b1, Mmax, temp_1} + {Mmin, temp_1}) ;
	
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

endmodule


//
// Description:	 Determine the normalization shift amount and perform 16-shift
//


module FPAddSub_NormalizeModule(
		Sum,
		Mmin,
		Shift
    );

	// Input ports
	input [`DWIDTH:0] Sum ;					// Mantissa sum including hidden 1 and GRS
	
	// Output ports
	output [`DWIDTH:0] Mmin ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount
	//Changes in this doesn't matter since even Bfloat16 can't go beyond 7 shift to the mantissa (only 3 bits valid here)  
	// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[16] ? 5'b00000 :	 
		Sum[15] ? 5'b00001 : 
		Sum[14] ? 5'b00010 : 
		Sum[13] ? 5'b00011 : 
		Sum[12] ? 5'b00100 : 
		Sum[11] ? 5'b00101 : 
		Sum[10] ? 5'b00110 : 
		Sum[9] ? 5'b00111 :
		Sum[8] ? 5'b01000 :
		Sum[7] ? 5'b01001 :
		Sum[6] ? 5'b01010 :
		Sum[5] ? 5'b01011 :
		Sum[4] ? 5'b01100 : 5'b01101
	//	Sum[19] ? 5'b01101 :
	//	Sum[18] ? 5'b01110 :
	//	Sum[17] ? 5'b01111 :
	//	Sum[16] ? 5'b10000 :
	//	Sum[15] ? 5'b10001 :
	//	Sum[14] ? 5'b10010 :
	//	Sum[13] ? 5'b10011 :
	//	Sum[12] ? 5'b10100 :
	//	Sum[11] ? 5'b10101 :
	//	Sum[10] ? 5'b10110 :
	//	Sum[9] ? 5'b10111 :
	//	Sum[8] ? 5'b11000 :
	//	Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [`DWIDTH:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[8:0], 8'b00000000} : Sum; 
	end
	
	// Assign outputs
	assign Mmin = Lvl1;						// Take out smaller mantissa

endmodule


// Description:	 Normalization shift stage 1, performs 12|8|4|3|2|1|0 shift
//
//Hardcoding loop start and end values of i. To avoid ODIN limitations. i=`DWIDTH*2+1 wasn't working.

module FPAddSub_NormalizeShift1(
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	input [`DWIDTH:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [3:0] Shift ;						// Shift amount
	
	// Output ports
	output [`DWIDTH:0] Mmin ;						// The smaller mantissa
	
	reg	  [`DWIDTH:0]		Lvl2;
	wire    [2*`DWIDTH+1:0]    Stage1;	
	reg	  [`DWIDTH:0]		Lvl3;
	wire    [2*`DWIDTH+1:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {MminP, MminP};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: Lvl2 <= Stage1[`DWIDTH:0];       		
			// Rotate by 4
			2'b01: begin for (i=33; i>=17; i=i-1) begin Lvl2[i-`DWIDTH -1] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
			// Rotate by 8
			2'b10: begin for (i=33; i>=17; i=i-1) begin Lvl2[i-`DWIDTH -1] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
			// Rotate by 12
			2'b11: begin for (i=33; i>=17; i=i-1) begin Lvl2[i-`DWIDTH -1] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[`DWIDTH:0];
			// Rotate by 1
			2'b01: begin for (i=33; i>=17; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
			// Rotate by 2
			2'b10: begin for (i=33; i>=17; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
			// Rotate by 3
			2'b11: begin for (i=33; i>=17; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
	  endcase
	end
	
	// Assign outputs
	assign Mmin = Lvl3;						// Take out smaller mantissa			
	
endmodule


// Description:	 Normalization shift stage 2, calculates post-normalization
//						 mantissa and exponent, as well as the bits used in rounding		
//


module FPAddSub_NormalizeShift2(
		PSSum,
		CExp,
		Shift,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [`DWIDTH:0] PSSum ;					// The Pre-Shift-Sum
	input [`EXPONENT-1:0] CExp ;
	input [4:0] Shift ;					// Amount to be shifted

	// Output ports
	output [`MANTISSA-1:0] NormM ;				// Normalized mantissa
	output [`EXPONENT:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;

	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [`EXPONENT:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [`EXPONENT:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = PSSum[`DWIDTH] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|PSSum ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[`EXPONENT] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = PSSum[`DWIDTH-1:`EXPONENT+1] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = PSSum[`EXPONENT] ; 
	assign R = PSSum[`EXPONENT-1] ;
	assign S = |PSSum[`EXPONENT-2:0] ;
	
endmodule


// Description:	 Performs 'Round to nearest, tie to even'-rounding on the
//						 normalized mantissa according to the G, R, S bits. Calculates
//						 final result and checks for exponent overflow.
//


module FPAddSub_RoundModule(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		Z,
		EOF
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [`EXPONENT:0] NormE ;				// Normalized exponent
	input [`MANTISSA-1:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	
	// Output ports
	output [`DWIDTH-1:0] Z ;					// Final result
	output EOF ;
	
	// Internal signals
	wire [`MANTISSA:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [`MANTISSA-1:0] RoundM ;				// The final rounded sum
	wire [`EXPONENT:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
        wire FSgn;
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	
	wire [`EXPONENT:0]temp_2;
	assign temp_2 = 0;
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[`MANTISSA-1:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[`MANTISSA] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? temp_2 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[`EXPONENT-1:0], RoundM[`MANTISSA-1:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[`EXPONENT];
	
endmodule


//
// Description:	 Check the final result for exception conditions and set
//						 flags accordingly.
//


module FPAddSub_ExceptionModule(
		Z,
		NegE,
		R,
		S,
		InputExc,
		EOF,
		P,
		Flags
    );
	 
	// Input ports
	input [`DWIDTH-1:0] Z	;					// Final product
	input NegE ;						// Negative exponent?
	input R ;							// Round bit
	input S ;							// Sticky bit
	input [4:0] InputExc ;			// Exceptions in inputs A and B
	input EOF ;
	
	// Output ports
	output [`DWIDTH-1:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[`MANTISSA+`EXPONENT-1:`MANTISSA]) & ~|(Z[`MANTISSA+`EXPONENT-1:`MANTISSA]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule
